magic
tech sky130A
magscale 1 2
timestamp 1698855384
<< error_p >>
rect 291918 364661 292030 364662
rect 291918 364581 292030 364582
<< metal3 >>
rect 511820 700416 514320 704810
rect 521432 700416 523932 703946
rect 511820 697916 523932 700416
rect 514086 669710 519258 697916
rect 134328 664538 519258 669710
rect 5373 337581 128286 337911
rect 344 337472 128286 337581
rect 5373 336821 128286 337472
rect 2990 294360 109888 295024
rect 342 294248 109888 294360
rect 2990 293144 109888 294248
rect 106790 282948 109888 293144
rect 6645 280718 102170 281808
rect 127196 280822 128286 336821
rect 6645 251338 7735 280718
rect 101936 280716 102170 280718
rect 342 251226 7735 251338
rect 6645 251087 7735 251226
rect 31331 277997 103188 279087
rect 31331 124117 32421 277997
rect 3945 123716 32421 124117
rect 326 123604 32421 123716
rect 3945 123027 32421 123604
rect 61553 275530 102104 276620
rect 61553 80603 62643 275530
rect 134328 274476 139500 664538
rect 572176 406600 582975 406686
rect 572176 406488 583606 406600
rect 572176 406300 582975 406488
rect 572176 374237 572562 406300
rect 1853 80494 62643 80603
rect 342 80382 62643 80494
rect 1853 79513 62643 80382
rect 74033 273716 102558 274146
rect 1115 37272 4017 37406
rect 342 37245 4017 37272
rect 74033 37245 74463 273716
rect 342 37160 74463 37245
rect 1115 36815 74463 37160
rect 87083 270683 102092 271773
rect 1115 36682 4017 36815
rect 87083 16181 88173 270683
rect 127280 269304 139500 274476
rect 154704 373851 572562 374237
rect 106618 236639 109716 266324
rect 115987 257334 116373 267445
rect 154704 257334 155090 373851
rect 115987 256948 155090 257334
rect 162337 364696 578379 366371
rect 162337 364661 581142 364696
rect 162337 364582 291918 364661
rect 292030 364584 581142 364661
rect 292030 364582 578379 364584
rect 162337 363273 578379 364582
rect 162337 236639 165435 363273
rect 291918 351954 292030 363273
rect 581030 360178 581142 364584
rect 581030 360066 583606 360178
rect 106618 233541 165435 236639
rect 1455 15850 88173 16181
rect 342 15738 88173 15850
rect 1455 15091 88173 15738
use pmu_circuits_top_level  pmu_circuits_top_level_0
timestamp 1698839394
transform 1 0 133834 0 1 279467
box -31742 -14099 -5382 4428
use user_analog_project_wrapper_pmu  user_analog_project_wrapper_pmu_0
timestamp 1698800988
transform 1 0 -26 0 1 10
box -800 -800 584800 704800
<< end >>

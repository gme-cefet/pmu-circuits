magic
tech sky130A
magscale 1 2
timestamp 1695834725
<< nwell >>
rect -430 1995 11477 3558
rect -430 1875 3662 1995
rect 9764 1990 11477 1995
rect -414 169 3662 1875
rect 9558 1617 11271 1626
rect 9558 85 11272 1617
<< psubdiff >>
rect -179 -270 -16 -219
rect 3226 -270 3405 -219
rect -179 -276 -91 -270
rect -179 -1052 -91 -951
rect 3317 -292 3405 -270
rect 3317 -1052 3405 -967
rect -179 -1121 -81 -1052
rect 3345 -1121 3405 -1052
<< nsubdiff >>
rect -394 3488 -334 3522
rect 11381 3488 11441 3522
rect -394 3462 -360 3488
rect -394 2065 -360 2091
rect 11407 3462 11441 3488
rect 11407 2065 11441 2091
rect -394 2031 -334 2065
rect 11381 2031 11441 2065
rect -378 1805 -318 1839
rect 3566 1805 3626 1839
rect -378 1779 -344 1805
rect -378 239 -344 265
rect 3592 1779 3626 1805
rect 3592 239 3626 265
rect -378 205 -318 239
rect 3566 205 3626 239
rect 9594 1547 9654 1581
rect 11176 1547 11236 1581
rect 9594 1521 9628 1547
rect 9594 155 9628 181
rect 11202 1521 11236 1547
rect 11202 155 11236 181
rect 9594 121 9654 155
rect 11176 121 11236 155
<< psubdiffcont >>
rect -16 -270 3226 -219
rect -179 -951 -91 -276
rect 3317 -967 3405 -292
rect -81 -1121 3345 -1052
<< nsubdiffcont >>
rect -334 3488 11381 3522
rect -394 2091 -360 3462
rect 11407 2091 11441 3462
rect -334 2031 11381 2065
rect -318 1805 3566 1839
rect -378 265 -344 1779
rect 3592 265 3626 1779
rect -318 205 3566 239
rect 9654 1547 11176 1581
rect 9594 181 9628 1521
rect 11202 181 11236 1521
rect 9654 121 11176 155
<< locali >>
rect -394 3488 -334 3522
rect 11381 3488 11441 3522
rect -394 3462 -360 3488
rect -360 3330 -199 3376
rect 369 3361 494 3488
rect 1153 3361 1278 3488
rect 1937 3361 2062 3488
rect 2721 3361 2846 3488
rect 3505 3361 3630 3488
rect 4289 3361 4414 3488
rect 5079 3358 5204 3488
rect 5863 3360 5988 3488
rect 6655 3362 6780 3488
rect 7439 3362 7564 3488
rect 8223 3362 8348 3488
rect 9007 3362 9132 3488
rect 9791 3362 9916 3488
rect 10575 3362 10700 3488
rect 11407 3462 11441 3488
rect 11269 3330 11407 3376
rect -360 2884 -199 2930
rect 4299 2798 4406 2895
rect 4299 2742 4320 2798
rect 4384 2742 4406 2798
rect -360 2630 -199 2676
rect 4299 2662 4406 2742
rect 5100 2816 5207 2893
rect 5874 2816 5981 2897
rect 5100 2720 5981 2816
rect 5100 2660 5207 2720
rect 5874 2664 5981 2720
rect 6660 2801 6767 2895
rect 11269 2884 11407 2930
rect 6660 2745 6682 2801
rect 6746 2745 6767 2801
rect 6660 2662 6767 2745
rect 11269 2630 11407 2676
rect -360 2184 -199 2230
rect 11269 2184 11407 2230
rect -394 2065 -360 2091
rect 11407 2065 11441 2091
rect -394 2031 -334 2065
rect 11381 2031 11441 2065
rect -374 1950 11423 2031
rect -325 1839 -47 1950
rect -378 1805 -318 1839
rect 3566 1805 3626 1839
rect -378 1779 -344 1805
rect -344 1634 2 1680
rect 385 1665 510 1805
rect 1175 1662 1300 1805
rect 1959 1664 2084 1805
rect 2751 1666 2876 1805
rect 3592 1779 3626 1805
rect 3260 1634 3592 1680
rect -344 1234 -243 1634
rect 3521 1234 3592 1634
rect -344 1188 2 1234
rect 395 1102 502 1199
rect 395 1046 416 1102
rect 480 1046 502 1102
rect -344 934 2 980
rect 395 966 502 1046
rect 1196 1120 1303 1197
rect 1970 1120 2077 1201
rect 1196 1024 2077 1120
rect 1196 964 1303 1024
rect 1970 968 2077 1024
rect 2756 1105 2863 1199
rect 3260 1188 3592 1234
rect 2756 1049 2778 1105
rect 2842 1049 2863 1105
rect 2756 966 2863 1049
rect 3260 946 3337 980
rect 3445 946 3592 980
rect 3260 934 3592 946
rect -344 534 -252 934
rect 3522 534 3592 934
rect -344 488 2 534
rect 124 442 158 534
rect 752 442 786 534
rect 124 408 786 442
rect 2476 426 2510 534
rect 3104 426 3138 534
rect 3260 522 3592 534
rect 3260 488 3337 522
rect 3445 488 3592 522
rect 2476 404 3284 426
rect 2476 392 3074 404
rect 3055 315 3074 392
rect 3254 315 3284 404
rect 3055 297 3284 315
rect -378 239 -344 265
rect 10384 1581 10616 1950
rect 3592 239 3626 265
rect -378 205 -318 239
rect 3566 205 3626 239
rect 9594 1547 9654 1581
rect 11176 1547 11236 1581
rect 9594 1521 9628 1547
rect 9763 1449 11055 1547
rect 11202 1521 11236 1547
rect 9594 155 9628 181
rect 11202 155 11236 181
rect 9594 121 9654 155
rect 11176 121 11236 155
rect -179 -276 -91 -260
rect -32 -270 -16 -219
rect 3226 -270 3242 -219
rect -450 -951 -179 -300
rect 3317 -292 3405 -276
rect -91 -429 317 -357
rect 452 -361 2732 -325
rect 2902 -429 3317 -357
rect 282 -937 317 -429
rect -91 -951 317 -937
rect -450 -964 317 -951
rect -180 -1009 317 -964
rect 282 -1052 317 -1009
rect 698 -1052 733 -429
rect 1114 -1052 1149 -429
rect 1530 -1052 1565 -429
rect 1946 -1052 1981 -429
rect 2362 -1052 2397 -429
rect 2778 -1052 2813 -429
rect 3194 -937 3229 -429
rect 2902 -967 3317 -937
rect 2902 -1009 3405 -967
rect 3194 -1052 3229 -1009
rect -97 -1121 -81 -1052
rect 3345 -1121 3361 -1052
<< viali >>
rect 4320 2742 4384 2798
rect 6682 2745 6746 2801
rect 416 1046 480 1102
rect 2778 1049 2842 1105
rect 3074 315 3254 404
<< metal1 >>
rect 776 2934 886 3326
rect 1554 2934 1676 3326
rect 2338 2934 2460 3326
rect 3122 2934 3244 3326
rect 3906 2934 4028 3326
rect 4690 2934 4812 3326
rect 5474 2934 5596 3326
rect 6258 2934 6380 3326
rect 7042 2934 7164 3326
rect 7826 2934 7948 3326
rect 8610 2934 8732 3326
rect 9394 2934 9516 3326
rect 10178 3258 10300 3326
rect 10178 3022 10192 3258
rect 10284 3022 10300 3258
rect 10178 2934 10300 3022
rect 373 2806 500 2891
rect 1157 2806 1284 2891
rect 1941 2806 2068 2891
rect 2725 2806 2852 2891
rect 3509 2806 3636 2891
rect 373 2801 3636 2806
rect 373 2746 3346 2801
rect 3628 2746 3636 2801
rect 373 2741 3636 2746
rect 373 2671 500 2741
rect 1157 2671 1284 2741
rect 1941 2671 2068 2741
rect 2725 2671 2852 2741
rect 3509 2671 3636 2741
rect 4299 2809 4406 2895
rect 6660 2809 6767 2895
rect 4299 2801 6767 2809
rect 4299 2798 6682 2801
rect 4299 2742 4320 2798
rect 4384 2745 6682 2798
rect 6746 2745 6767 2801
rect 4384 2742 6767 2745
rect 4299 2731 6767 2742
rect 4299 2662 4406 2731
rect 6660 2662 6767 2731
rect 7429 2806 7556 2889
rect 8213 2806 8340 2889
rect 8997 2806 9124 2889
rect 9781 2806 9908 2889
rect 10565 2806 10692 2889
rect 7429 2801 10692 2806
rect 7429 2746 7437 2801
rect 7719 2746 10692 2801
rect 7429 2741 10692 2746
rect 7429 2669 7556 2741
rect 8213 2669 8340 2741
rect 8997 2669 9124 2741
rect 9781 2669 9908 2741
rect 10565 2669 10692 2741
rect 64 1963 124 2627
rect 776 2234 886 2626
rect 1554 2234 1676 2626
rect 2338 2234 2460 2626
rect 3122 2234 3244 2626
rect 3906 2234 4028 2626
rect 4690 2234 4812 2626
rect 5474 2234 5596 2626
rect 6258 2234 6380 2626
rect 7042 2234 7164 2626
rect 7826 2234 7948 2626
rect 8610 2234 8732 2626
rect 9394 2234 9516 2626
rect 10178 2234 10300 2626
rect 189 2154 3825 2178
rect 189 2135 1056 2154
rect 973 2102 1056 2135
rect 2968 2135 3825 2154
rect 2968 2102 3041 2135
rect 973 2082 3041 2102
rect 4290 1995 4397 2199
rect 4893 2131 6177 2178
rect 5482 1995 5587 2131
rect 64 1895 3755 1963
rect 4289 1956 4398 1995
rect -471 1736 3144 1768
rect -471 399 -406 1736
rect 118 1630 164 1736
rect 746 1630 792 1736
rect 902 1630 948 1736
rect 1530 1630 1576 1736
rect 1686 1630 1732 1736
rect 2314 1630 2360 1736
rect 2470 1630 2516 1736
rect 3098 1630 3144 1736
rect 395 1113 502 1199
rect 2756 1113 2863 1199
rect 395 1105 2863 1113
rect 395 1102 2778 1105
rect 395 1046 416 1102
rect 480 1049 2778 1102
rect 2842 1049 2863 1105
rect 480 1046 2863 1049
rect 395 1035 2863 1046
rect 395 966 502 1035
rect 2756 966 2863 1035
rect 792 538 902 930
rect 1576 538 1686 930
rect 2360 538 2470 930
rect 386 399 493 503
rect 989 422 2273 482
rect 2752 430 2859 505
rect -471 382 493 399
rect -471 347 301 382
rect -464 346 301 347
rect 266 299 301 346
rect 461 348 493 382
rect 461 299 492 348
rect 266 285 492 299
rect 1546 -15 1693 422
rect 2753 397 2859 430
rect 3055 404 3284 426
rect 2635 379 2861 397
rect 2635 296 2668 379
rect 2828 296 2861 379
rect 3055 315 3074 404
rect 3254 391 3284 404
rect 3687 391 3755 1895
rect 4171 1936 4513 1956
rect 4171 1846 4233 1936
rect 4453 1846 4513 1936
rect 4171 1825 4513 1846
rect 5481 1742 5587 1995
rect 6656 1958 6763 2201
rect 7245 2154 10881 2178
rect 7245 2135 8112 2154
rect 8029 2102 8112 2135
rect 10024 2135 10881 2154
rect 10024 2102 10097 2135
rect 8029 2082 10097 2102
rect 6656 1957 6800 1958
rect 6573 1937 6915 1957
rect 6573 1847 6635 1937
rect 6855 1847 6915 1937
rect 6573 1826 6915 1847
rect 10967 1913 11011 2625
rect 10967 1844 11439 1913
rect 10354 951 10464 1399
rect 9767 808 11051 951
rect 9767 755 10267 808
rect 10551 755 11051 808
rect 3254 321 3755 391
rect 3254 315 3284 321
rect 3055 297 3284 315
rect 10354 307 10464 699
rect 11324 315 11439 1844
rect 11095 307 11444 315
rect 2635 283 2861 296
rect 9680 251 9767 307
rect 10267 251 10551 307
rect 11051 253 11444 307
rect 11051 251 11446 253
rect 9680 214 11446 251
rect 9680 208 11138 214
rect 770 -88 2068 -15
rect 40 -1011 236 -965
rect 365 -1119 418 -433
rect 770 -933 820 -88
rect 1345 -203 1721 -172
rect 1345 -304 1413 -203
rect 1661 -304 1721 -203
rect 1345 -309 1721 -304
rect 1186 -355 1896 -309
rect 1186 -933 1236 -355
rect 1602 -933 1652 -355
rect 2018 -933 2068 -88
rect 2432 -234 3543 -171
rect 2434 -933 2484 -234
rect 3444 -875 3543 -234
rect 11260 -736 11446 214
rect 11126 -793 11474 -736
rect 3439 -907 3699 -875
rect 452 -1011 2732 -965
rect 2948 -1011 3144 -965
rect 3439 -1119 3473 -907
rect 365 -1172 3473 -1119
rect 3670 -1172 3699 -907
rect 365 -1184 3699 -1172
rect 397 -1185 3699 -1184
rect 3439 -1197 3699 -1185
rect 11126 -1143 11187 -793
rect 11424 -1143 11474 -793
rect 11126 -1199 11474 -1143
<< via1 >>
rect 10192 3022 10284 3258
rect 3346 2746 3628 2801
rect 7437 2746 7719 2801
rect 1056 2102 2968 2154
rect 301 299 461 382
rect 2668 296 2828 379
rect 4233 1846 4453 1936
rect 8112 2102 10024 2154
rect 6635 1847 6855 1937
rect 1413 -304 1661 -203
rect 3473 -1172 3670 -907
rect 11187 -1143 11424 -793
<< metal2 >>
rect 10138 3258 10340 3326
rect 10138 3022 10192 3258
rect 10284 3022 10340 3258
rect 10138 2934 10340 3022
rect 3338 2801 7727 2806
rect 3338 2746 3346 2801
rect 3628 2746 7437 2801
rect 7719 2746 7727 2801
rect 3338 2741 7727 2746
rect 10187 2172 10282 2934
rect 973 2154 10282 2172
rect 973 2102 1056 2154
rect 2968 2102 8112 2154
rect 10024 2102 10282 2154
rect 973 2082 10282 2102
rect 6573 1957 6915 1958
rect 3779 1937 6915 1957
rect 3779 1936 6635 1937
rect 3779 1846 4233 1936
rect 4453 1847 6635 1936
rect 6855 1847 6915 1937
rect 4453 1846 6915 1847
rect 3779 1828 6915 1846
rect 3779 1827 6773 1828
rect 266 382 492 399
rect 266 299 301 382
rect 461 378 492 382
rect 2635 379 2861 397
rect 2635 378 2668 379
rect 461 303 2668 378
rect 461 299 492 303
rect 266 285 492 299
rect 2635 296 2668 303
rect 2828 296 2861 379
rect 2635 283 2861 296
rect 3779 130 3881 1827
rect 8132 1787 8442 2082
rect 2152 20 3881 130
rect 1345 -181 1721 -172
rect 2154 -181 2248 20
rect 3779 19 3881 20
rect 1345 -203 2248 -181
rect 1345 -304 1413 -203
rect 1661 -258 2248 -203
rect 1661 -304 1721 -258
rect 1345 -322 1721 -304
rect 11126 -793 11474 -736
rect 3439 -907 3699 -875
rect 3439 -1172 3473 -907
rect 3670 -1054 3699 -907
rect 11126 -1054 11187 -793
rect 3670 -1143 11187 -1054
rect 11424 -1143 11474 -793
rect 3670 -1172 11474 -1143
rect 3439 -1197 11474 -1172
rect 3477 -1198 11474 -1197
rect 11126 -1199 11474 -1198
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_8
timestamp 1695788690
transform 1 0 3048 0 1 -683
box -158 -338 158 338
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_9
timestamp 1695788690
transform 1 0 2216 0 1 -683
box -158 -338 158 338
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_10
timestamp 1695788690
transform 1 0 2632 0 1 -683
box -158 -338 158 338
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_11
timestamp 1695788690
transform 1 0 1384 0 1 -683
box -158 -338 158 338
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_12
timestamp 1695788690
transform 1 0 1800 0 1 -683
box -158 -338 158 338
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_13
timestamp 1695788690
transform 1 0 552 0 1 -683
box -158 -338 158 338
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_14
timestamp 1695788690
transform 1 0 968 0 1 -683
box -158 -338 158 338
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_15
timestamp 1695788690
transform 1 0 136 0 1 -683
box -158 -338 158 338
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_0
timestamp 1695405779
transform 0 1 455 -1 0 734
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_1
timestamp 1695405779
transform 0 1 1239 -1 0 734
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_2
timestamp 1695405779
transform 0 1 2023 -1 0 734
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_3
timestamp 1695405779
transform 0 1 2807 -1 0 734
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_4
timestamp 1695405779
transform 0 1 455 -1 0 1434
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_5
timestamp 1695405779
transform 0 1 1239 -1 0 1434
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_6
timestamp 1695405779
transform 0 1 2023 -1 0 1434
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_7
timestamp 1695405779
transform 0 1 2807 -1 0 1434
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_8
timestamp 1695405779
transform 0 1 3575 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_9
timestamp 1695405779
transform 0 1 2791 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_10
timestamp 1695405779
transform 0 1 5143 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_11
timestamp 1695405779
transform 0 1 4359 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_12
timestamp 1695405779
transform 0 1 3575 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_13
timestamp 1695405779
transform 0 1 2791 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_14
timestamp 1695405779
transform 0 1 5143 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_15
timestamp 1695405779
transform 0 1 4359 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_16
timestamp 1695405779
transform 0 1 1223 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_17
timestamp 1695405779
transform 0 1 1223 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_18
timestamp 1695405779
transform 0 1 2007 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_19
timestamp 1695405779
transform 0 1 2007 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_20
timestamp 1695405779
transform 0 1 5927 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_21
timestamp 1695405779
transform 0 1 6711 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_22
timestamp 1695405779
transform 0 1 5927 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_23
timestamp 1695405779
transform 0 1 6711 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_26
timestamp 1695405779
transform 0 1 7495 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_27
timestamp 1695405779
transform 0 1 7495 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_30
timestamp 1695405779
transform 0 1 9847 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_31
timestamp 1695405779
transform 0 1 9847 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_32
timestamp 1695405779
transform 0 1 439 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_33
timestamp 1695405779
transform 0 1 439 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_34
timestamp 1695405779
transform 0 1 10631 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_35
timestamp 1695405779
transform 0 1 10631 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_36
timestamp 1695405779
transform 0 1 9063 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_37
timestamp 1695405779
transform 0 1 9063 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_38
timestamp 1695405779
transform 0 1 8279 -1 0 2430
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_39
timestamp 1695405779
transform 0 1 8279 -1 0 3130
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_40
timestamp 1695405779
transform 0 1 10017 -1 0 503
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_41
timestamp 1695405779
transform 0 1 10801 -1 0 503
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_42
timestamp 1695405779
transform 0 1 10017 -1 0 1203
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_NTRJ8S  sky130_fd_pr__pfet_01v8_lvt_NTRJ8S_43
timestamp 1695405779
transform 0 1 10801 -1 0 1203
box -294 -350 294 350
use sky130_fd_pr__pfet_01v8_lvt_WCVK8S  sky130_fd_pr__pfet_01v8_lvt_WCVK8S_0
timestamp 1695405779
transform 0 1 3391 -1 0 734
box -294 -150 294 150
use sky130_fd_pr__pfet_01v8_lvt_WCVK8S  sky130_fd_pr__pfet_01v8_lvt_WCVK8S_1
timestamp 1695405779
transform 0 1 3391 -1 0 1434
box -294 -150 294 150
use sky130_fd_pr__pfet_01v8_lvt_WCVK8S  sky130_fd_pr__pfet_01v8_lvt_WCVK8S_2
timestamp 1695405779
transform 0 -1 -129 -1 0 1434
box -294 -150 294 150
use sky130_fd_pr__pfet_01v8_lvt_WCVK8S  sky130_fd_pr__pfet_01v8_lvt_WCVK8S_3
timestamp 1695405779
transform 0 -1 -129 -1 0 734
box -294 -150 294 150
use sky130_fd_pr__pfet_01v8_lvt_WCVK8S  sky130_fd_pr__pfet_01v8_lvt_WCVK8S_4
timestamp 1695405779
transform 0 -1 -145 -1 0 2430
box -294 -150 294 150
use sky130_fd_pr__pfet_01v8_lvt_WCVK8S  sky130_fd_pr__pfet_01v8_lvt_WCVK8S_5
timestamp 1695405779
transform 0 -1 -145 -1 0 3130
box -294 -150 294 150
use sky130_fd_pr__pfet_01v8_lvt_WCVK8S  sky130_fd_pr__pfet_01v8_lvt_WCVK8S_6
timestamp 1695405779
transform 0 1 11215 -1 0 2430
box -294 -150 294 150
use sky130_fd_pr__pfet_01v8_lvt_WCVK8S  sky130_fd_pr__pfet_01v8_lvt_WCVK8S_7
timestamp 1695405779
transform 0 1 11215 -1 0 3130
box -294 -150 294 150
<< labels >>
rlabel metal2 8173 1828 8383 1963 3 Ip2
rlabel metal1 5502 1758 5575 1808 3 Iref
rlabel metal1 1575 -10 1648 40 3 Vg
rlabel metal2 355 304 428 354 3 Ip1
rlabel locali -360 -740 -255 -614 3 SS
rlabel locali 10477 1727 10551 1815 3 DD
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1697036621
<< error_p >>
rect 2598 1528 2644 1540
rect 2598 1468 2604 1528
rect 2638 1468 2644 1528
rect 2598 1230 2644 1242
rect 2598 1170 2604 1230
rect 2638 1170 2644 1230
rect 2454 294 2536 298
<< nwell >>
rect 2885 169 3563 1835
<< psubdiff >>
rect -230 1743 -206 1833
rect 2708 1743 2732 1833
rect 2701 402 2819 426
rect 2701 260 2819 284
<< nsubdiff >>
rect 2921 1765 2981 1799
rect 3467 1765 3527 1799
rect 2921 1739 2955 1765
rect 2921 239 2955 265
rect 3493 1739 3527 1765
rect 3493 239 3527 265
rect 2921 205 2981 239
rect 3467 205 3527 239
<< psubdiffcont >>
rect -206 1743 2708 1833
rect 2701 284 2819 402
<< nsubdiffcont >>
rect 2981 1765 3467 1799
rect 2921 265 2955 1739
rect 3493 265 3527 1739
rect 2981 205 3467 239
<< locali >>
rect 2448 1833 2732 1838
rect -222 1743 -206 1833
rect 2708 1743 2732 1833
rect 2448 1738 2732 1743
rect 2921 1765 2981 1799
rect 3467 1765 3527 1799
rect 2921 1739 2955 1765
rect -200 1634 1094 1670
rect -200 1310 -158 1634
rect 1460 1590 2921 1636
rect 1298 1422 1338 1450
rect 1298 1382 1682 1422
rect -14 1346 1246 1382
rect -200 1274 1094 1310
rect -200 950 -158 1274
rect 1210 1042 1246 1346
rect 1298 1128 1338 1382
rect 2700 1332 2740 1590
rect 1460 1286 2740 1332
rect 2790 1275 2862 1299
rect 2790 1192 2808 1275
rect 2843 1192 2862 1275
rect 1298 1086 1730 1128
rect 2790 1061 2862 1192
rect 2358 1042 2862 1061
rect 1210 1025 2862 1042
rect 1210 1022 2540 1025
rect -14 1008 2540 1022
rect -14 986 1298 1008
rect -200 914 1094 950
rect -200 590 -158 914
rect 1238 662 1298 986
rect 1432 684 2712 718
rect -14 626 1298 662
rect 1238 620 1298 626
rect -200 554 1094 590
rect 1238 586 2540 620
rect 1238 302 1280 586
rect -14 266 1280 302
rect 2676 418 2712 684
rect 2676 402 2819 418
rect 2676 298 2701 402
rect 2536 294 2701 298
rect 1432 284 2701 294
rect 1432 269 2819 284
rect 1502 268 2819 269
rect 1502 264 2712 268
rect 3396 1739 3527 1765
rect 3396 1681 3493 1739
rect 3004 1333 3042 1619
rect 3404 1377 3441 1619
rect 3270 1355 3457 1377
rect 3004 1294 3175 1333
rect 3119 1238 3175 1294
rect 3270 1307 3334 1355
rect 3431 1307 3457 1355
rect 3270 1292 3457 1307
rect 3271 1238 3327 1292
rect 3042 941 3076 1051
rect 3370 964 3404 1051
rect 3331 942 3436 964
rect 3331 941 3351 942
rect 3042 893 3351 941
rect 3042 765 3076 893
rect 3331 874 3351 893
rect 3414 874 3436 942
rect 3331 857 3436 874
rect 3370 765 3404 857
rect 1502 125 2488 264
rect 2921 239 2955 265
rect 3118 239 3328 354
rect 3493 239 3527 265
rect 2921 205 2981 239
rect 3467 205 3527 239
<< viali >>
rect 2476 1751 2703 1820
rect 2808 1192 2843 1275
rect 3334 1307 3431 1355
rect 3351 874 3414 942
<< metal1 >>
rect 2448 1837 2732 1838
rect 2448 1820 3249 1837
rect 2448 1751 2476 1820
rect 2703 1751 3249 1820
rect 2448 1748 3249 1751
rect 2448 1738 2732 1748
rect 1185 1674 1390 1716
rect 510 1638 2861 1674
rect 3190 1647 3249 1748
rect 1340 1634 2861 1638
rect -130 352 -88 1584
rect 1168 866 1210 1584
rect 1340 1378 1388 1634
rect 2793 1605 2861 1634
rect 2793 1545 3061 1605
rect 2793 1544 2861 1545
rect 2644 1378 2692 1540
rect 1340 1334 2692 1378
rect 3203 1352 3247 1430
rect 1340 1170 1388 1334
rect 2644 1170 2692 1334
rect 2790 1307 3247 1352
rect 3309 1359 3496 1377
rect 3309 1307 3334 1359
rect 3432 1307 3496 1359
rect 2790 1275 2862 1307
rect 3309 1292 3496 1307
rect 2790 1192 2808 1275
rect 2843 1192 2862 1275
rect 2790 1176 2862 1192
rect 2309 1084 2809 1125
rect 2774 969 2809 1084
rect 3186 969 3256 1007
rect 1316 866 1358 960
rect 1168 804 1358 866
rect 1168 756 1210 804
rect 1168 536 1212 756
rect 1316 674 1358 804
rect 2614 674 2656 960
rect 2774 885 3256 969
rect 3186 800 3256 885
rect 3331 942 3436 964
rect 3331 874 3351 942
rect 3414 874 3436 942
rect 3331 857 3436 874
rect 1316 636 2656 674
rect 1168 482 1210 536
rect 1316 482 1358 636
rect 1168 420 1358 482
rect 1168 352 1210 420
rect 1316 344 1358 420
rect 2614 543 2656 636
rect 2614 486 3052 543
rect 2614 410 3048 486
rect 2614 344 2656 410
<< via1 >>
rect 3334 1355 3432 1359
rect 3334 1307 3431 1355
rect 3431 1307 3432 1355
rect 3351 874 3414 942
<< metal2 >>
rect 3309 1363 3496 1377
rect 3309 1307 3334 1363
rect 3437 1307 3496 1363
rect 3309 1292 3496 1307
rect 3331 942 3436 964
rect 3331 874 3351 942
rect 3414 874 3436 942
rect 3331 857 3436 874
<< via2 >>
rect 3334 1359 3437 1363
rect 3334 1307 3432 1359
rect 3432 1307 3437 1359
rect 3351 874 3414 942
<< metal3 >>
rect 3309 1363 3496 1377
rect 3309 1307 3334 1363
rect 3437 1307 3496 1363
rect 3309 1292 3496 1307
rect 3307 942 3460 990
rect 3307 874 3351 942
rect 3414 874 3460 942
rect 3307 839 3460 874
use sky130_fd_pr__nfet_01v8_lvt_62AYNZ  sky130_fd_pr__nfet_01v8_lvt_62AYNZ_0
timestamp 1695672277
transform 0 1 1986 -1 0 864
box -158 -638 158 638
use sky130_fd_pr__nfet_01v8_lvt_62AYNZ  sky130_fd_pr__nfet_01v8_lvt_62AYNZ_1
timestamp 1695672277
transform 0 1 1986 -1 0 440
box -158 -638 158 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_4
timestamp 1697035654
transform 0 -1 540 1 0 1508
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_5
timestamp 1697035654
transform 0 -1 540 1 0 1148
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_6
timestamp 1697035654
transform 0 -1 540 1 0 788
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_7
timestamp 1697035654
transform 0 -1 540 1 0 428
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P34KHJ  sky130_fd_pr__nfet_01v8_lvt_P34KHJ_0
timestamp 1695675331
transform 0 -1 2016 -1 0 1206
box -98 -638 98 638
use sky130_fd_pr__nfet_01v8_lvt_P34KHJ  sky130_fd_pr__nfet_01v8_lvt_P34KHJ_1
timestamp 1695675331
transform 0 -1 2016 -1 0 1504
box -98 -638 98 638
use sky130_fd_pr__pfet_01v8_lvt_G2G9KE  sky130_fd_pr__pfet_01v8_lvt_G2G9KE_0
timestamp 1697034391
transform 0 -1 3223 1 0 1131
box -174 -200 174 200
use sky130_fd_pr__pfet_01v8_lvt_G2G9KE  sky130_fd_pr__pfet_01v8_lvt_G2G9KE_1
timestamp 1697034391
transform 0 -1 3223 1 0 1539
box -174 -200 174 200
use sky130_fd_pr__pfet_01v8_lvt_NCVK88  sky130_fd_pr__pfet_01v8_lvt_NCVK88_0
timestamp 1695678748
transform 0 1 3223 -1 0 565
box -294 -200 294 200
<< labels >>
rlabel metal1 2763 429 2838 493 3 IN
rlabel locali 1811 1758 1886 1822 3 SS
rlabel locali 3425 1704 3463 1738 3 DD
rlabel metal1 1248 1664 1292 1703 3 OUT
<< end >>

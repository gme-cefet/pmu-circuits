magic
tech sky130A
timestamp 1696460965
<< end >>

* NGSPICE file created from ldo.ext - technology: sky130A

.subckt ldo DD SS Iref VB VS OUT
X0 a_9110_n8196.t1 VB a_8766_n8196.t0 SS sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=5.19 l=1.43
X1 SS Iref a_9110_n8196.t7 SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X2 DD.t17 a_8766_n8196.t4 OUT.t4 DD.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.9 as=1.5 ps=10.9 w=5.17 l=0.37
X3 DD.t9 DD.t6 DD.t8 DD.t7 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.258 ps=2.36 w=0.89 l=3.89
X4 a_9110_n8196.t6 Iref SS SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X5 a_8766_n8196.t5 OUT.t3 sky130_fd_pr__cap_mim_m3_1 l=15 w=4
X6 DD.t1 a_9330_n9998.t4 a_9330_n9998.t5 DD.t0 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X7 DD.t13 a_9330_n9998.t6 a_8766_n8196.t3 DD.t12 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X8 SS Iref a_9330_n9998.t1 SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X9 SS SS SS SS sky130_fd_pr__nfet_01v8_lvt ad=17.7 pd=129 as=1.48 ps=10.8 w=5.1 l=0.66
X10 OUT.t2 VS a_9110_n8196.t2 OUT.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.76 pd=12.7 as=1.76 ps=12.7 w=6.07 l=1.27
X11 a_9110_n8196.t5 Iref SS SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X12 SS Iref Iref SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X13 DD.t11 a_9330_n9998.t7 a_8766_n8196.t2 DD.t10 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X14 OUT.t1 VS a_9110_n8196.t3 OUT.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.76 pd=12.7 as=1.76 ps=12.7 w=6.07 l=1.27
X15 SS Iref a_9110_n8196.t4 SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X16 a_9110_n8196.t0 VB a_8766_n8196.t1 SS sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=5.19 l=1.43
X17 DD.t5 DD.t2 DD.t4 DD.t3 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0 ps=0 w=0.89 l=3.89
X18 SS SS SS SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=0 ps=0 w=5.1 l=0.66
X19 DD.t15 a_9330_n9998.t2 a_9330_n9998.t3 DD.t14 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X20 a_9330_n9998.t0 Iref SS SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X21 Iref Iref SS SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
R0 a_8766_n8196.n0 a_8766_n8196.t4 191.636
R1 a_8766_n8196.n0 a_8766_n8196.t2 34.661
R2 a_8766_n8196.n0 a_8766_n8196.t3 33.291
R3 a_8766_n8196.t0 a_8766_n8196.n2 4.51459
R4 a_8766_n8196.n2 a_8766_n8196.t1 3.35375
R5 a_8766_n8196.n1 a_8766_n8196.n0 2.51069
R6 a_8766_n8196.n2 a_8766_n8196.n1 1.37236
R7 a_8766_n8196.n1 a_8766_n8196.t5 0.251842
R8 a_9110_n8196.n0 a_9110_n8196.t2 7.40825
R9 a_9110_n8196.n0 a_9110_n8196.t3 4.70699
R10 a_9110_n8196.n1 a_9110_n8196.t4 4.53569
R11 a_9110_n8196.n4 a_9110_n8196.t5 4.53369
R12 a_9110_n8196.t6 a_9110_n8196.n5 4.38957
R13 a_9110_n8196.n2 a_9110_n8196.t7 4.3873
R14 a_9110_n8196.n3 a_9110_n8196.t0 4.26166
R15 a_9110_n8196.n3 a_9110_n8196.t1 4.06962
R16 a_9110_n8196.n5 a_9110_n8196.n2 2.26478
R17 a_9110_n8196.n4 a_9110_n8196.n3 2.0915
R18 a_9110_n8196.n1 a_9110_n8196.n0 0.66715
R19 a_9110_n8196.n5 a_9110_n8196.n4 0.1505
R20 a_9110_n8196.n2 a_9110_n8196.n1 0.144506
R21 OUT.n1 OUT.n2 336.49
R22 OUT.n0 OUT.t1 7.2144
R23 OUT.n3 OUT.t4 5.74557
R24 OUT.n0 OUT.t2 4.7068
R25 OUT.n1 OUT.t0 4.25837
R26 OUT.n3 OUT.t3 0.292821
R27 OUT.n3 OUT.n1 0.234051
R28 OUT OUT.n3 0.221825
R29 OUT.n1 OUT.n0 0.0894987
R30 DD.n2 DD.n6 459.673
R31 DD.t3 DD.t12 367.363
R32 DD.t0 DD.t10 367.363
R33 DD.n3 DD.n0 254.948
R34 DD.n1 DD.t3 232.912
R35 DD.n0 DD.t7 213.075
R36 DD.n2 DD.t0 193.233
R37 DD.n10 DD.n9 186.632
R38 DD.n2 DD.t14 174.131
R39 DD.n12 DD.t16 73.8353
R40 DD.n11 DD.t5 60.0995
R41 DD.n6 DD.t9 60.0995
R42 DD.n12 DD.n11 53.4946
R43 DD.n3 DD.t8 48.3828
R44 DD.n9 DD.t4 45.276
R45 DD.n5 DD.n4 34.174
R46 DD.n8 DD.n7 34.174
R47 DD.n8 DD.t13 32.0995
R48 DD.n7 DD.t15 32.0995
R49 DD.n5 DD.t1 32.0995
R50 DD.n4 DD.t11 32.0995
R51 DD.n4 DD.n3 28.5054
R52 DD.n9 DD.n8 28.5054
R53 DD.n2 DD.n5 18.0327
R54 DD.n7 DD.n2 16.1447
R55 DD.n0 DD.t6 9.484
R56 DD.n1 DD.t2 9.47999
R57 DD.n13 DD.n12 8.40959
R58 DD.n14 DD.n10 8.10924
R59 DD.t16 DD.t17 5.52608
R60 DD.n14 DD.n13 5.40633
R61 DD.n10 DD.n1 0.844913
R62 DD DD.n14 0.190885
R63 a_9330_n9998.n1 a_9330_n9998.t5 32.4466
R64 a_9330_n9998.n0 a_9330_n9998.t3 32.4466
R65 a_9330_n9998.t4 a_9330_n9998.t7 19.1411
R66 a_9330_n9998.t2 a_9330_n9998.t6 19.1411
R67 a_9330_n9998.t1 a_9330_n9998.n4 10.1828
R68 a_9330_n9998.n3 a_9330_n9998.t4 9.48031
R69 a_9330_n9998.n2 a_9330_n9998.t2 9.48031
R70 a_9330_n9998.n4 a_9330_n9998.n1 5.92365
R71 a_9330_n9998.n4 a_9330_n9998.t0 5.36911
R72 a_9330_n9998.n0 a_9330_n9998.n2 0.351043
R73 a_9330_n9998.n1 a_9330_n9998.n3 0.351043
R74 a_9330_n9998.n1 a_9330_n9998.n0 0.100294
C0 Iref OUT 0.0248f
C1 Iref VS 0.00227f
C2 OUT VB 1.47f
C3 VB VS 0.134f
C4 DD OUT 1.35f
C5 DD VS 0.00151f
C6 Iref VB 0.267f
C7 OUT VS 2.28f
C8 DD VB 0.0106f
C9 Iref SS 8.14f
C10 VS SS 0.71f
C11 VB SS 4.08f
C12 OUT SS 11.8f
C13 DD SS 20.7f
C14 a_9330_n9998.n0 SS 0.0865f
C15 a_9330_n9998.n1 SS 0.923f
C16 a_9330_n9998.t0 SS 0.159f
C17 a_9330_n9998.t6 SS 0.706f
C18 a_9330_n9998.t2 SS 0.421f
C19 a_9330_n9998.n2 SS 0.225f
C20 a_9330_n9998.t3 SS 0.00544f
C21 a_9330_n9998.t7 SS 0.706f
C22 a_9330_n9998.t4 SS 0.421f
C23 a_9330_n9998.n3 SS 0.225f
C24 a_9330_n9998.t5 SS 0.00544f
C25 a_9330_n9998.n4 SS 1.07f
C26 a_9330_n9998.t1 SS 0.344f
C27 DD.n0 SS 0.336f
C28 DD.n1 SS 0.312f
C29 DD.t16 SS 0.633f
C30 DD.n2 SS 0.335f
C31 DD.t6 SS 0.161f
C32 DD.t7 SS 0.31f
C33 DD.t8 SS 0.00749f
C34 DD.n3 SS 0.0477f
C35 DD.t11 SS 0.00157f
C36 DD.n4 SS 0.0623f
C37 DD.t1 SS 0.00157f
C38 DD.n5 SS 0.0544f
C39 DD.t14 SS 0.289f
C40 DD.t10 SS 0.392f
C41 DD.t0 SS 0.299f
C42 DD.t9 SS 0.00741f
C43 DD.n6 SS 0.0317f
C44 DD.t15 SS 0.00157f
C45 DD.n7 SS 0.053f
C46 DD.t13 SS 0.00157f
C47 DD.n8 SS 0.0623f
C48 DD.t4 SS 0.00469f
C49 DD.n9 SS 0.0471f
C50 DD.t2 SS 0.161f
C51 DD.t12 SS 0.392f
C52 DD.t3 SS 0.32f
C53 DD.n10 SS 0.212f
C54 DD.t17 SS 0.00909f
C55 DD.t5 SS 0.00741f
C56 DD.n11 SS 0.0289f
C57 DD.n12 SS 0.204f
C58 DD.n13 SS 0.0791f
C59 DD.n14 SS 0.292f
C60 OUT.n0 SS 0.357f
C61 OUT.n1 SS 2.66f
C62 OUT.t4 SS 0.0208f
C63 OUT.t3 SS 5.29f
C64 OUT.t0 SS 0.0439f
C65 OUT.t1 SS 0.133f
C66 OUT.t2 SS 0.0215f
C67 OUT.n2 SS 0.674f
C68 OUT.n3 SS 0.396f
C69 a_9110_n8196.t7 SS 0.0644f
C70 a_9110_n8196.t4 SS 0.0716f
C71 a_9110_n8196.t2 SS 0.144f
C72 a_9110_n8196.t3 SS 0.0219f
C73 a_9110_n8196.n0 SS 0.546f
C74 a_9110_n8196.n1 SS 0.418f
C75 a_9110_n8196.n2 SS 0.243f
C76 a_9110_n8196.t0 SS 0.0908f
C77 a_9110_n8196.t1 SS 0.0757f
C78 a_9110_n8196.n3 SS 0.875f
C79 a_9110_n8196.t5 SS 0.0714f
C80 a_9110_n8196.n4 SS 0.471f
C81 a_9110_n8196.n5 SS 0.243f
C82 a_9110_n8196.t6 SS 0.0645f
C83 a_8766_n8196.n0 SS 0.631f
C84 a_8766_n8196.t4 SS 0.0546f
C85 a_8766_n8196.t2 SS 0.00656f
C86 a_8766_n8196.t3 SS 0.00418f
C87 a_8766_n8196.t5 SS 5.2f
C88 a_8766_n8196.n1 SS 0.901f
C89 a_8766_n8196.t1 SS 0.0181f
C90 a_8766_n8196.n2 SS 0.704f
C91 a_8766_n8196.t0 SS 0.0787f
.ends


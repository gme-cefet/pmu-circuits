magic
tech sky130A
magscale 1 2
timestamp 1698328096
<< psubdiff >>
rect -3409 39 -3339 205
rect 8950 39 9048 205
rect -3409 -111 -3256 39
rect 8895 -84 9048 39
rect 3980 -2357 4095 -1928
rect 3980 -4178 4095 -4154
rect -3256 -5028 -3127 -4904
rect 8739 -5005 8895 -4904
rect 8739 -5028 9048 -5005
rect 8895 -5029 9048 -5028
rect -3409 -5056 -3256 -5032
<< psubdiffcont >>
rect -3339 39 8950 205
rect -3409 -5032 -3256 -111
rect 3980 -4154 4095 -2357
rect -3127 -5028 8739 -4904
rect 8895 -5005 9048 -84
<< locali >>
rect -3409 39 -3339 205
rect 8950 39 9048 205
rect -3409 -111 -3256 39
rect 8895 -84 9048 39
rect -3123 -164 8690 -108
rect -3171 -252 8690 -164
rect -3171 -1646 -3003 -252
rect 8596 -1413 8673 -252
rect 8428 -1570 8673 -1413
rect -2486 -1626 -2093 -1611
rect -957 -1626 -564 -1603
rect -147 -1626 246 -1607
rect -3179 -1681 -3003 -1646
rect -2839 -1634 755 -1626
rect 837 -1634 940 -1630
rect -3179 -3407 -3051 -1681
rect -2839 -1797 940 -1634
rect -2839 -1800 755 -1797
rect 837 -3395 940 -1797
rect 6753 -1644 6871 -1640
rect 6753 -1650 7072 -1644
rect 6753 -1706 7766 -1650
rect 1428 -1965 1589 -1919
rect 2237 -1965 2445 -1917
rect 1428 -2007 2445 -1965
rect 1428 -2058 2409 -2007
rect 1469 -2110 2409 -2058
rect 3921 -2357 4108 -1879
rect 6753 -2048 7158 -1706
rect 7834 -1817 8683 -1570
rect 6753 -2057 7766 -2048
rect 6753 -2117 6871 -2057
rect 7054 -2088 7766 -2057
rect 5090 -2231 6356 -2118
rect 6501 -2177 6871 -2117
rect 6501 -2178 6857 -2177
rect 3921 -2409 3980 -2357
rect 2371 -2649 2445 -2587
rect 3023 -3102 3314 -3070
rect 3023 -3283 3056 -3102
rect 3269 -3103 3314 -3102
rect 3269 -3278 3529 -3103
rect 3269 -3283 3314 -3278
rect 3023 -3314 3314 -3283
rect -3256 -3853 1471 -3684
rect -3256 -3886 -2777 -3853
rect 497 -3859 1444 -3853
rect 497 -3886 1468 -3859
rect -3256 -3965 -2836 -3886
rect 572 -3960 1468 -3886
rect -3256 -4581 -3131 -3965
rect 634 -4136 1468 -3960
rect 4095 -2409 4108 -2357
rect 6481 -2344 6869 -2178
rect 6481 -2364 6873 -2344
rect 6483 -3175 6873 -2364
rect 6501 -3215 6857 -3175
rect 4095 -4148 4625 -4030
rect 3980 -4170 4095 -4154
rect -3014 -4904 -2449 -4567
rect 463 -4904 653 -4604
rect 1428 -4614 1604 -4467
rect 1612 -4614 2191 -4489
rect 1428 -4616 2208 -4614
rect 2236 -4616 2383 -4583
rect 1428 -4904 2438 -4616
rect 4265 -4904 4625 -4148
rect -3256 -5028 -3127 -4904
rect 8739 -5005 8895 -4904
rect 8739 -5028 9048 -5005
rect 8891 -5029 9048 -5028
rect -3409 -5048 -3256 -5032
<< viali >>
rect 7158 -2048 7770 -1706
rect 3056 -3283 3269 -3102
<< metal1 >>
rect 2619 -2211 2953 -1472
rect 7108 -1706 7820 -1654
rect 7108 -2048 7158 -1706
rect 7770 -2048 7820 -1706
rect 7108 -2092 7820 -2048
rect 2619 -2248 3216 -2211
rect 2619 -2413 2666 -2248
rect 3172 -2413 3216 -2248
rect 2619 -2444 3216 -2413
rect 1203 -2899 1271 -2875
rect -34 -3452 77 -3270
rect 1203 -3452 1303 -2899
rect 3023 -3102 3314 -3070
rect 3023 -3283 3056 -3102
rect 3269 -3283 3314 -3102
rect 3023 -3314 3314 -3283
rect -34 -3546 1303 -3452
rect -712 -3699 993 -3631
rect 907 -4253 993 -3699
rect 3114 -3989 3219 -3314
rect 2795 -4072 3219 -3989
rect 2799 -4175 3219 -4072
rect 907 -4319 1360 -4253
rect 1282 -4778 1360 -4319
<< via1 >>
rect 7158 -2048 7770 -1706
rect 2666 -2413 3172 -2248
<< metal2 >>
rect 8493 -1604 9031 189
rect 8492 -1626 9031 -1604
rect 7108 -1706 7820 -1654
rect 5386 -1934 5601 -1765
rect 1273 -2026 5601 -1934
rect 1273 -2048 5600 -2026
rect 7108 -2048 7158 -1706
rect 7770 -1756 7820 -1706
rect 8492 -1756 9032 -1626
rect 7770 -1966 9032 -1756
rect 7770 -2048 7820 -1966
rect 1273 -2495 1349 -2048
rect 7108 -2092 7820 -2048
rect 2589 -2240 3269 -2183
rect 2589 -2575 2663 -2240
rect 3202 -2575 3269 -2240
rect 2589 -2614 3269 -2575
<< via2 >>
rect 2663 -2248 3202 -2240
rect 2663 -2413 2666 -2248
rect 2666 -2413 3172 -2248
rect 3172 -2413 3202 -2248
rect 2663 -2575 3202 -2413
<< metal3 >>
rect 2589 -2240 3269 -2183
rect 2589 -2575 2663 -2240
rect 3202 -2575 3269 -2240
rect 2589 -2614 3269 -2575
rect 2973 -4749 3260 -2614
rect 6759 -4404 8187 -3699
rect 5770 -4588 8187 -4404
rect 5770 -4749 6048 -4588
rect 2973 -4943 6048 -4749
use iref_2nA_igenerator  iref_2nA_igenerator_0
timestamp 1695828444
transform 0 -1 -101 -1 0 1852
box 3769 -3056 6630 -1355
use iref_2nA_mirrors  iref_2nA_mirrors_0
timestamp 1695834725
transform 1 0 -2745 0 1 -3616
box -471 -1199 11477 3558
use iref_2nA_vref  iref_2nA_vref_0
timestamp 1697059543
transform -1 0 5067 0 1 -1039
box -1459 -3811 1752 -845
<< labels >>
flabel metal2 8592 -558 8796 -328 0 FreeSans 1600 0 0 0 DD
port 0 nsew
flabel metal3 7304 -4258 7508 -4028 0 FreeSans 1600 0 0 0 IREF
port 1 nsew
flabel locali -3140 -3898 -2976 -3750 0 FreeSans 1600 0 0 0 SS
port 2 nsew
<< end >>

magic
tech sky130A
timestamp 1696344833
<< nmoslvt >>
rect -33 -255 33 255
<< ndiff >>
rect -62 249 -33 255
rect -62 -249 -56 249
rect -39 -249 -33 249
rect -62 -255 -33 -249
rect 33 249 62 255
rect 33 -249 39 249
rect 56 -249 62 249
rect 33 -255 62 -249
<< ndiffc >>
rect -56 -249 -39 249
rect 39 -249 56 249
<< poly >>
rect -33 291 33 299
rect -33 274 -25 291
rect 25 274 33 291
rect -33 255 33 274
rect -33 -274 33 -255
rect -33 -291 -25 -274
rect 25 -291 33 -274
rect -33 -299 33 -291
<< polycont >>
rect -25 274 25 291
rect -25 -291 25 -274
<< locali >>
rect -33 274 -25 291
rect 25 274 33 291
rect -56 249 -39 257
rect -56 -257 -39 -249
rect 39 249 56 257
rect 39 -257 56 -249
rect -33 -291 -25 -274
rect 25 -291 33 -274
<< viali >>
rect -25 274 25 291
rect -56 -249 -39 249
rect 39 -249 56 249
rect -25 -291 25 -274
<< metal1 >>
rect -31 291 31 294
rect -31 274 -25 291
rect 25 274 31 291
rect -31 271 31 274
rect -59 249 -36 255
rect -59 -249 -56 249
rect -39 -249 -36 249
rect -59 -255 -36 -249
rect 36 249 59 255
rect 36 -249 39 249
rect 56 -249 59 249
rect 36 -255 59 -249
rect -31 -274 31 -271
rect -31 -291 -25 -274
rect 25 -291 31 -274
rect -31 -294 31 -291
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.10 l 0.66 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

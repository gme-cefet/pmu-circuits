magic
tech sky130A
magscale 1 2
timestamp 1695345667
<< nwell >>
rect -532 -337 532 337
<< pmos >>
rect -438 -237 438 237
<< pdiff >>
rect -496 225 -438 237
rect -496 -225 -484 225
rect -450 -225 -438 225
rect -496 -237 -438 -225
rect 438 225 496 237
rect 438 -225 450 225
rect 484 -225 496 225
rect 438 -237 496 -225
<< pdiffc >>
rect -484 -225 -450 225
rect 450 -225 484 225
<< poly >>
rect -438 318 438 334
rect -438 284 -422 318
rect 422 284 438 318
rect -438 237 438 284
rect -438 -284 438 -237
rect -438 -318 -422 -284
rect 422 -318 438 -284
rect -438 -334 438 -318
<< polycont >>
rect -422 284 422 318
rect -422 -318 422 -284
<< locali >>
rect -438 284 -422 318
rect 422 284 438 318
rect -484 225 -450 241
rect -484 -241 -450 -225
rect 450 225 484 241
rect 450 -241 484 -225
rect -438 -318 -422 -284
rect 422 -318 438 -284
<< viali >>
rect -422 284 422 318
rect -484 -225 -450 225
rect 450 -225 484 225
rect -422 -318 422 -284
<< metal1 >>
rect -434 318 434 324
rect -434 284 -422 318
rect 422 284 434 318
rect -434 278 434 284
rect -490 225 -444 237
rect -490 -225 -484 225
rect -450 -225 -444 225
rect -490 -237 -444 -225
rect 444 225 490 237
rect 444 -225 450 225
rect 484 -225 490 225
rect 444 -237 490 -225
rect -434 -284 434 -278
rect -434 -318 -422 -284
rect 422 -318 434 -284
rect -434 -324 434 -318
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.37 l 4.38 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1698839394
<< locali >>
rect -8382 -4309 -5382 -3944
rect -8382 -11125 -8044 -4309
rect -5779 -11125 -5382 -4309
rect -8382 -11445 -5382 -11125
<< viali >>
rect -8044 -11125 -5779 -4309
<< metal1 >>
rect -28038 4206 -20162 4428
rect -28038 2956 -27694 4206
rect -20419 2956 -20162 4206
rect -28038 2784 -20162 2956
rect -31736 2187 -30575 2343
rect -31736 1380 -31586 2187
rect -30717 1807 -30575 2187
rect -30717 1628 -27982 1807
rect -30717 1380 -30575 1628
rect -31736 1253 -30575 1380
rect -29735 -1290 -27800 -1085
rect -31736 -2989 -30575 -2846
rect -31736 -3786 -31573 -2989
rect -30742 -3258 -30575 -2989
rect -29735 -3258 -29530 -1290
rect -30742 -3463 -29530 -3258
rect -28980 -2070 -27480 -1641
rect -30742 -3786 -30575 -3463
rect -31736 -3936 -30575 -3786
rect -31277 -5322 -29518 -5321
rect -28980 -5322 -28551 -2070
rect -31277 -5397 -28551 -5322
rect -31277 -5695 -31213 -5397
rect -28630 -5695 -28551 -5397
rect -31277 -5751 -28551 -5695
rect -8382 -4309 -5382 -3944
rect -8382 -11125 -8044 -4309
rect -5779 -11125 -5382 -4309
rect -22861 -12701 -22275 -11251
rect -8382 -11445 -5382 -11125
rect -29548 -12906 -22247 -12701
rect -29548 -13943 -29355 -12906
rect -22499 -13943 -22247 -12906
rect -29548 -14099 -22247 -13943
<< via1 >>
rect -27694 2956 -20419 4206
rect -31586 1380 -30717 2187
rect -31573 -3786 -30742 -2989
rect -31213 -5695 -28630 -5397
rect -8044 -11125 -5779 -4309
rect -29355 -13943 -22499 -12906
<< metal2 >>
rect -28038 4206 -20162 4428
rect -28038 2956 -27694 4206
rect -20419 2956 -20162 4206
rect -28038 2784 -20162 2956
rect -31736 2187 -30575 2343
rect -31736 1380 -31586 2187
rect -30717 1380 -30575 2187
rect -31736 1253 -30575 1380
rect -31736 -2989 -30575 -2846
rect -31736 -3786 -31573 -2989
rect -30742 -3786 -30575 -2989
rect -31736 -3936 -30575 -3786
rect -8382 -4309 -5382 -3944
rect -31277 -5397 -28551 -5322
rect -31277 -5695 -31213 -5397
rect -28630 -5695 -28551 -5397
rect -31277 -5751 -28551 -5695
rect -29147 -7013 -26556 -6782
rect -31742 -7860 -30581 -7694
rect -31742 -8645 -31579 -7860
rect -30764 -8020 -30581 -7860
rect -29147 -8020 -28916 -7013
rect -30764 -8251 -28916 -8020
rect -30764 -8645 -30581 -8251
rect -31742 -8784 -30581 -8645
rect -8382 -11125 -8044 -4309
rect -5779 -11125 -5382 -4309
rect -8382 -11445 -5382 -11125
rect -21636 -11954 -21456 -11483
rect -21636 -12004 -16976 -11954
rect -21636 -12106 -21591 -12004
rect -17029 -12106 -16976 -12004
rect -21636 -12134 -16976 -12106
rect -29548 -12906 -22247 -12701
rect -29548 -13943 -29355 -12906
rect -22499 -13943 -22247 -12906
rect -29548 -14099 -22247 -13943
<< via2 >>
rect -27694 2956 -20419 4206
rect -31586 1380 -30717 2187
rect -31573 -3786 -30742 -2989
rect -31213 -5695 -28630 -5397
rect -31579 -8645 -30764 -7860
rect -8044 -11125 -5779 -4309
rect -21591 -12106 -17029 -12004
rect -29355 -13943 -22499 -12906
<< metal3 >>
rect -28038 4206 -20162 4428
rect -28038 2956 -27694 4206
rect -20419 2956 -20162 4206
rect -28038 2784 -20162 2956
rect -31736 2187 -30575 2343
rect -31736 1380 -31586 2187
rect -30717 1380 -30575 2187
rect -31736 1253 -30575 1380
rect -6638 1355 -5477 2445
rect -6586 501 -5835 1355
rect -31248 -201 -27862 30
rect -31248 -380 -31017 -201
rect -9200 -250 -5835 501
rect -31736 -1470 -30575 -380
rect -31736 -2989 -30575 -2846
rect -31736 -3786 -31573 -2989
rect -30742 -3786 -30575 -2989
rect -31736 -3936 -30575 -3786
rect -8382 -4309 -5382 -3944
rect -31277 -5397 -28551 -5322
rect -31277 -5695 -31213 -5397
rect -28630 -5695 -28551 -5397
rect -31277 -5751 -28551 -5695
rect -31742 -7860 -30581 -7694
rect -31742 -8645 -31579 -7860
rect -30764 -8645 -30581 -7860
rect -31742 -8784 -30581 -8645
rect -8382 -11125 -8044 -4309
rect -5779 -11125 -5382 -4309
rect -8382 -11445 -5382 -11125
rect -21636 -12004 -16976 -11954
rect -21636 -12106 -21591 -12004
rect -17029 -12106 -16976 -12004
rect -21636 -12134 -16976 -12106
rect -29548 -12906 -22247 -12701
rect -29548 -13943 -29355 -12906
rect -22499 -13943 -22247 -12906
rect -29548 -14099 -22247 -13943
use pmu_circuits  pmu_circuits_0
timestamp 1698332589
transform -1 0 -9223 0 -1 8924
box -1074 5482 18938 20761
<< end >>

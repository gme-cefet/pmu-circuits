magic
tech sky130A
magscale 1 2
timestamp 1697065484
<< nwell >>
rect 4896 -5413 4913 2917
<< psubdiff >>
rect 3945 3035 5864 3126
rect 848 2887 1106 2915
rect 1002 2825 1106 2887
rect 3945 2820 4068 3035
rect 5741 2820 5864 3035
rect 8694 2887 8961 2915
rect 8694 2825 8807 2887
rect 1002 1159 1126 1249
rect 8694 1159 8807 1249
rect 1002 -507 1127 -417
rect 8694 -507 8807 -417
rect 1002 -2173 1128 -2083
rect 8694 -2173 8807 -2083
rect 1002 -3839 1106 -3749
rect 8694 -3839 8807 -3749
rect 1002 -5521 1131 -5513
rect 848 -5593 1131 -5521
rect 8773 -5521 8807 -5513
rect 8773 -5593 8961 -5521
<< psubdiffcont >>
rect 848 -5521 1002 2887
rect 1131 -5593 8773 -5513
rect 8807 -5521 8961 2887
<< locali >>
rect 848 2887 1002 2903
rect 1253 2868 3484 3386
rect 4732 3169 5079 3214
rect 4732 2793 4779 3169
rect 5025 2793 5079 3169
rect 8694 2825 8695 2915
rect 8807 2887 8961 2903
rect 4732 2761 5079 2793
rect 4863 -5377 4946 2761
rect 8694 1159 8695 1249
rect 8694 -507 8695 -417
rect 8694 -2173 8695 -2083
rect 8694 -3839 8695 -3749
rect 2838 -5513 3824 -5444
rect 5985 -5513 6971 -5451
rect 1002 -5521 1131 -5513
rect 848 -5593 1131 -5521
rect 8773 -5521 8807 -5513
rect 8773 -5593 8961 -5521
<< viali >>
rect 4779 2793 5025 3169
<< metal1 >>
rect 5904 3283 6208 3583
rect 4869 3277 8080 3283
rect 4732 3169 8080 3277
rect 4732 2793 4779 3169
rect 5025 3046 8080 3169
rect 5025 2793 5079 3046
rect 4732 2761 5079 2793
<< metal2 >>
rect 4448 2984 4574 3823
rect 4109 2941 4574 2984
rect 4108 2927 4574 2941
rect 4108 2479 4248 2927
rect 4108 2365 4798 2479
rect 5016 2458 5683 2459
rect 5016 2374 5704 2458
rect 4751 1954 5059 2032
rect 5600 375 5704 2374
rect 4107 282 4772 367
rect 5037 290 5704 375
rect 4107 -873 4219 282
rect 4107 -958 4793 -873
rect 5016 -874 5683 -873
rect 5016 -958 5704 -874
rect 5600 -2957 5704 -958
rect 4107 -3046 4772 -2961
rect 5037 -3042 5704 -2957
rect 4107 -4205 4219 -3046
rect 4107 -4290 4793 -4205
rect 5016 -4290 5685 -4205
rect 4760 -4679 4938 -4627
rect 4858 -5421 4938 -4679
rect 5594 -5421 5685 -4290
rect 4858 -5485 5685 -5421
<< metal3 >>
rect 4105 1951 4772 2036
rect 4105 794 4217 1951
rect 4105 709 4793 794
rect 5016 792 5683 793
rect 5016 708 5704 792
rect 5600 -1291 5704 708
rect 4104 -1386 4769 -1301
rect 5037 -1376 5704 -1291
rect 4104 -2539 4216 -1386
rect 4104 -2624 4793 -2539
rect 5016 -2540 5683 -2539
rect 5016 -2624 5704 -2540
rect 5600 -4623 5704 -2624
rect 5037 -4708 5704 -4623
use mdls_inv  mdls_inv_0
timestamp 1697036621
transform -1 0 8473 0 1 -5582
box -230 125 3563 1838
use mdls_inv  mdls_inv_1
timestamp 1697036621
transform 1 0 1336 0 1 -5582
box -230 125 3563 1838
use mdls_inv  mdls_inv_2
timestamp 1697036621
transform -1 0 8473 0 1 1082
box -230 125 3563 1838
use mdls_inv  mdls_inv_3
timestamp 1697036621
transform 1 0 1336 0 1 1082
box -230 125 3563 1838
use mdls_inv  mdls_inv_4
timestamp 1697036621
transform 1 0 1336 0 1 -584
box -230 125 3563 1838
use mdls_inv  mdls_inv_5
timestamp 1697036621
transform -1 0 8473 0 1 -584
box -230 125 3563 1838
use mdls_inv  mdls_inv_6
timestamp 1697036621
transform 1 0 1336 0 1 -2250
box -230 125 3563 1838
use mdls_inv  mdls_inv_7
timestamp 1697036621
transform -1 0 8473 0 1 -2250
box -230 125 3563 1838
use mdls_inv  mdls_inv_8
timestamp 1697036621
transform 1 0 1336 0 1 -3916
box -230 125 3563 1838
use mdls_inv  mdls_inv_9
timestamp 1697036621
transform -1 0 8473 0 1 -3916
box -230 125 3563 1838
use ring_100mV_buffer  ring_100mV_buffer_0
timestamp 1697038384
transform 1 0 -2319 0 1 7075
box 3175 -3762 10387 -140
<< labels >>
flabel locali 1652 2982 2000 3234 0 FreeSans 1600 0 0 0 SS
port 0 nsew
flabel metal1 6454 3092 6660 3282 0 FreeSans 1600 0 0 0 DD
port 1 nsew
flabel space 7086 4956 7292 5146 0 FreeSans 1600 0 0 0 OUT
port 2 nsew
<< end >>

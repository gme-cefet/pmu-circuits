magic
tech sky130A
magscale 1 2
timestamp 1698861079
<< metal3 >>
rect 572176 406600 582975 406686
rect 572176 406488 583606 406600
rect 572176 406300 582975 406488
rect 572176 374237 572562 406300
rect 154704 373851 572562 374237
rect 5373 337581 128286 337911
rect 344 337472 128286 337581
rect 5373 336821 128286 337472
rect 2990 294360 109888 295024
rect 342 294248 109888 294360
rect 2990 293144 109888 294248
rect 106790 282948 109888 293144
rect 6645 280718 102170 281808
rect 127196 280822 128286 336821
rect 6645 251338 7735 280718
rect 101936 280716 102170 280718
rect 342 251226 7735 251338
rect 6645 251087 7735 251226
rect 31331 277997 103188 279087
rect 31331 124117 32421 277997
rect 3945 123716 32421 124117
rect 326 123604 32421 123716
rect 3945 123027 32421 123604
rect 61553 275530 102104 276620
rect 61553 80603 62643 275530
rect 134328 274476 139500 350418
rect 1853 80494 62643 80603
rect 342 80382 62643 80494
rect 1853 79513 62643 80382
rect 74033 273716 102558 274146
rect 1115 37272 4017 37406
rect 342 37245 4017 37272
rect 74033 37245 74463 273716
rect 342 37160 74463 37245
rect 1115 36815 74463 37160
rect 87083 270683 102092 271773
rect 1115 36682 4017 36815
rect 87083 16181 88173 270683
rect 127280 269304 139500 274476
rect 106618 236639 109716 266324
rect 115987 257334 116373 267445
rect 154704 257334 155090 373851
rect 115987 256948 155090 257334
rect 162337 364696 578379 366371
rect 162337 364584 581142 364696
rect 162337 363273 578379 364584
rect 162337 236639 165435 363273
rect 581030 360178 581142 364584
rect 581030 360066 583606 360178
rect 106618 233541 165435 236639
rect 1455 15850 88173 16181
rect 342 15738 88173 15850
rect 1455 15091 88173 15738
use pmu_circuits_top_level  pmu_circuits_top_level_0
timestamp 1698839394
transform 1 0 133834 0 1 279467
box -31742 -14099 -5382 4428
<< labels >>
flabel metal3 10028 336906 11894 337768 0 FreeSans 8000 0 0 0 gpio_noesd[11]
port 0 nsew
flabel metal3 9412 293530 11278 294392 0 FreeSans 8000 0 0 0 gpio_noesd[12]
port 1 nsew
flabel metal3 6760 251254 7466 251912 0 FreeSans 8000 0 0 0 gpio_noesd[13]
port 2 nsew
flabel metal3 7748 123292 8454 123950 0 FreeSans 8000 0 0 0 gpio_noesd[14]
port 3 nsew
flabel metal3 7280 79630 7986 80288 0 FreeSans 8000 0 0 0 gpio_noesd[15]
port 4 nsew
flabel metal3 6896 36870 8062 37110 0 FreeSans 8000 0 0 0 gpio_noesd[16]
port 5 nsew
flabel metal3 6686 15490 7852 15730 0 FreeSans 8000 0 0 0 gpio_noesd[17]
port 6 nsew
flabel metal3 573308 364318 574122 364838 0 FreeSans 8000 0 0 0 gpio_noesd[2]
port 7 nsew
flabel metal3 575802 406322 576204 406584 0 FreeSans 8000 0 0 0 gpio_noesd[3]
port 8 nsew
flabel metal3 135612 346104 138678 348766 0 FreeSans 12800 0 0 0 vssa1
port 9 nsew
<< end >>

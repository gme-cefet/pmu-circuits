* NGSPICE file created from aux.ext - technology: sky130A

.subckt aux gpio_analog[0] gpio_analog[10] gpio_analog[11] gpio_analog[12] gpio_analog[13]
+ gpio_analog[14] gpio_analog[15] gpio_analog[16] gpio_analog[17] gpio_analog[1] gpio_analog[2]
+ gpio_analog[3] gpio_analog[4] gpio_analog[5] gpio_analog[6] gpio_analog[7] gpio_analog[8]
+ gpio_analog[9] gpio_noesd[0] gpio_noesd[10] gpio_noesd[11] gpio_noesd[12] gpio_noesd[13]
+ gpio_noesd[14] gpio_noesd[15] gpio_noesd[16] gpio_noesd[17] gpio_noesd[1] gpio_noesd[2]
+ gpio_noesd[3] gpio_noesd[4] gpio_noesd[5] gpio_noesd[6] gpio_noesd[7] gpio_noesd[8]
+ gpio_noesd[9] io_analog[0] io_analog[10] io_analog[1] io_analog[2] io_analog[3]
+ io_analog[7] io_analog[8] io_analog[9] io_analog[4] io_analog[5] io_analog[6] io_clamp_high[0]
+ io_clamp_high[1] io_clamp_high[2] io_clamp_low[0] io_clamp_low[1] io_clamp_low[2]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9]
+ io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12] io_in_3v3[13] io_in_3v3[14]
+ io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18] io_in_3v3[19] io_in_3v3[1]
+ io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23] io_in_3v3[24] io_in_3v3[25]
+ io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4] io_in_3v3[5] io_in_3v3[6] io_in_3v3[7]
+ io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[2] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[16] io_out[17] io_out[18] io_out[19]
+ io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26]
+ io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101]
+ la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108]
+ la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114]
+ la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120]
+ la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69]
+ la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81]
+ la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88]
+ la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94]
+ la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2
+ user_irq[0] user_irq[1] user_irq[2] vccd2 vdda2 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i vssa1 io_out[15] vccd1 vdda1
X0 vccd1.t57 a_337443_613718.t2 a_337443_613718.t3 vccd1.t55 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X1 a_339370_613888.t9 a_335807_622237.t6 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t8 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X2 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_343294_619079# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X3 vccd1.t66 a_350942_613328.t6 a_350378_615130.t3 vccd1.t65 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X4 a_337674_621712# a_335807_622237.t7 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t3 vccd1.t7 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X5 a_337443_613718.t1 a_335807_622237.t2 a_335807_622237.t3 vccd1.t50 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X6 a_339370_613888.t8 a_335807_622237.t8 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t4 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X7 a_343294_617413# pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t5 vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X8 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT vssa1 vssa1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
R0 io_oeb[15] vssd1 sky130_fd_pr__res_generic_m3 w=0.56 l=0.6
X9 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t5 a_341600_622217.t7 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
R1 io_analog[4] io_clamp_high[0] sky130_fd_pr__res_generic_m3 w=11 l=0.25
X10 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_345642_615404# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X11 gpio_analog[3].t15 a_341600_622217.t10 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X12 vdda1 a_341600_622217.t11 gpio_analog[3].t19 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X13 a_341818_614929.t1 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t5 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X14 a_339370_613888.t7 a_335807_622237.t9 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t3 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X15 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t3 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t6 a_341818_616595.t5 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X16 a_350722_615130.t7 gpio_analog[7].t4 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X17 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t4 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t5 a_341818_613263.t5 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X18 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t2 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t7 a_341818_616595.t4 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X19 a_343294_620745# pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X20 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT a_345642_618736# vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X21 vccd1.t68 a_350942_613328.t7 a_350378_615130.t2 vccd1.t67 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X22 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_345642_616040.t6 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X23 io_out[15].t2 io_out[16].t0 a_350722_615130.t0 io_out[15].t0 sky130_fd_pr__pfet_01v8_lvt ad=1.76 pd=12.7 as=1.76 ps=12.7 w=6.07 l=1.27
X24 io_out[11].t0 a_352038_622652.t4 a_352038_622652.t5 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.499 pd=4.02 as=0.499 ps=4.02 w=1.72 l=3.1
X25 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t3 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_341818_619927.t5 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X26 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=100 ps=733 w=2.5 l=1
X27 a_339370_618592# a_335807_622237.t10 io_out[11].t3 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X28 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t2 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_341818_619927.t4 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X29 a_345642_613738# pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X30 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_345642_616040.t5 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X31 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.725 ps=5.58 w=2.5 l=1
X32 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t6 a_341600_622217.t6 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X33 a_341818_613263.t1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t6 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X34 a_345642_617706.t5 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X35 gpio_analog[3].t14 a_341600_622217.t12 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X36 a_343294_619079# pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t5 vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X37 a_345642_617070# pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X38 gpio_analog[3].t13 a_341600_622217.t13 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X39 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg a_335719_622037.t6 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X40 a_345642_616040.t1 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X41 a_337443_613718.t0 a_335807_622237.t0 a_335807_622237.t1 vccd1.t50 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X42 a_339370_613888.t6 a_335807_622237.t11 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t2 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X43 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t6 a_341818_618261.t4 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X44 a_350722_615130.t6 gpio_analog[7].t5 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X45 vccd1.t59 a_352038_622652.t2 a_352038_622652.t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.89
X46 vccd1.t40 vccd1.t38 vccd1.t39 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=2
R2 vssd1 io_oeb[11] sky130_fd_pr__res_generic_m3 w=0.56 l=0.58
X47 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t7 a_341818_618261.t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X48 a_339370_613888.t5 a_335807_622237.t12 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t11 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X49 gpio_analog[3].t12 a_341600_622217.t14 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X50 gpio_analog[3].t18 a_341600_622217.t15 vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X51 a_345642_620402# pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X52 vccd1.t47 a_350942_613328.t2 a_350942_613328.t3 vccd1.t46 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X53 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_345642_617706.t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
R3 vssa1 io_clamp_low[1] sky130_fd_pr__res_generic_m3 w=11 l=0.25
X54 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t8 a_343294_615747# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X55 a_336843_616061.t1 w_336471_617254# pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT vccd1.t43 sky130_fd_pr__pfet_01v8_lvt ad=0.995 pd=7.44 as=0.995 ps=7.44 w=3.43 l=2.77
X56 gpio_analog[3].t11 a_341600_622217.t16 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X57 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t7 a_345642_613738# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X58 vccd1.t69 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t12 a_339370_613888.t19 vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X59 vssa1 gpio_analog[7].t6 a_350722_615130.t5 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X60 a_345642_618736# pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X61 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t6 a_343294_614081# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X62 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_345642_617706.t2 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X63 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_345642_617070# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X64 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg a_335719_622037.t7 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X65 a_341818_618261.t6 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t8 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X66 vccd1.t70 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t13 a_339370_613888.t18 vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X67 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT a_345642_620402# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X68 vccd1.t71 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t14 a_339370_613888.t17 vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X69 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t7 a_341600_622217.t5 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X70 gpio_analog[3].t10 a_341600_622217.t17 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X71 a_345642_621038.t1 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
R4 io_oeb[16] vssd1 sky130_fd_pr__res_generic_m3 w=0.56 l=0.31
X72 vccd1.t75 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t4 a_337674_622496# vccd1.t21 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X73 gpio_analog[3].t17 a_341600_622217.t18 vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X74 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t2 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t8 a_341818_613263.t4 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X75 vccd1.t51 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t15 a_339370_613888.t16 vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X76 gpio_analog[3].t9 a_341600_622217.t19 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X77 vssa1 gpio_analog[7].t2 gpio_analog[7].t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X78 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT a_345642_619372.t4 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
R5 vssa1 io_clamp_low[0] sky130_fd_pr__res_generic_m3 w=11 l=0.25
X79 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t9 a_341818_616595.t6 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X80 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t8 a_343294_620745# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X81 a_345642_614374.t2 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X82 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t3 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t9 a_341818_613263.t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X83 vccd1.t37 vccd1.t35 vccd1.t36 vccd1.t21 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=2
R6 vssd1 io_oeb[12] sky130_fd_pr__res_generic_m3 w=0.56 l=0.49
X84 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t10 a_341818_613263.t2 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X85 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_345642_617070# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X86 vssa1 a_352038_622652.t6 io_out[11].t1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.238 pd=2.22 as=0.238 ps=2.22 w=0.82 l=1.05
X87 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t9 a_341600_622217.t4 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X88 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_345642_618736# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X89 vccd1.t52 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t16 a_339370_618592# vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X90 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t1 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_341818_619927.t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X91 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t4 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t7 a_341818_614929.t5 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X92 gpio_analog[3].t8 a_341600_622217.t20 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X93 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_343294_619079# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X94 a_339370_613888.t4 a_335807_622237.t13 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t10 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X95 vccd1.t34 vccd1.t31 vccd1.t33 vccd1.t32 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0 ps=0 w=0.89 l=3.89
X96 a_343294_615747# pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t8 vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X97 a_341818_616595.t1 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t9 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X98 a_339370_613888.t3 a_335807_622237.t14 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t9 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X99 gpio_analog[7].t1 gpio_analog[7].t0 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X100 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t1 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t9 a_341818_614929.t4 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X101 vccd1.t53 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t17 a_339370_613888.t15 vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X102 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t10 a_341818_618261.t2 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X103 a_341818_614929.t0 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t10 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X104 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t0 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t11 a_341818_614929.t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X105 a_345642_621038.t0 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X106 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t2 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t12 a_343294_615747# vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X107 vccd1.t76 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t5 a_337674_622496# vccd1.t21 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X108 vccd1.t30 vccd1.t28 vccd1.t29 vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=2
X109 a_337674_622496# a_335807_622237.t15 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg vccd1.t7 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X110 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_345642_617706.t6 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X111 a_335807_622237.t4 a_335719_622037.t8 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X112 vccd1.t60 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t18 a_339370_613888.t14 vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X113 a_339370_617808# a_335807_622237.t16 a_335719_622037.t5 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
R7 vssa1 io_clamp_high[2] sky130_fd_pr__res_generic_m3 w=11 l=0.25
X114 gpio_analog[3].t7 a_341600_622217.t21 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X115 vssa1 gpio_analog[7].t7 a_350942_613328.t5 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X116 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_345642_617706.t1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X117 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t0 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_345642_614374.t6 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X118 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_345642_617706.t0 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X119 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0 ps=0 w=2.5 l=1
X120 a_345642_619372.t6 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X121 a_339370_617808# a_335807_622237.t17 a_335719_622037.t4 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X122 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_345642_621038.t5 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X123 vccd1.t19 vccd1.t17 vccd1.t18 vccd1.t7 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=2
X124 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_345642_621038.t4 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X125 a_345642_615404# pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X126 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t0 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_341818_619927.t2 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X127 gpio_analog[3].t6 a_341600_622217.t22 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X128 vccd1.t27 vccd1.t24 vccd1.t26 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=2
X129 a_339370_613888.t2 a_335807_622237.t18 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t7 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X130 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_345642_615404# vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X131 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t4 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t10 a_343294_617413# vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X132 a_339370_618592# a_335807_622237.t19 io_out[11].t2 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X133 a_339370_613888.t1 a_335807_622237.t20 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t6 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X134 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT a_345642_619372.t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X135 a_345642_617706.t4 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X136 a_341818_619927.t1 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X137 vssa1 gpio_analog[7].t8 a_350722_615130.t4 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X138 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_345642_615404# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X139 a_335719_622037.t3 a_335719_622037.t2 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X140 a_337674_622496# a_335807_622237.t21 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg vccd1.t7 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X141 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT a_345642_619372.t2 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X142 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg a_336716_619863# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X143 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t13 a_341818_613263.t6 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X144 vccd1.t23 vccd1.t20 vccd1.t22 vccd1.t21 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=2
X145 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t10 a_341600_622217.t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X146 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t11 a_345642_613738# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X147 gpio_analog[3].t5 a_341600_622217.t23 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X148 a_341818_613263.t0 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t12 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X149 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t11 a_341818_619927.t6 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X150 vccd1.t63 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t6 a_337674_621712# vccd1.t21 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X151 vccd1.t16 vccd1.t14 a_336843_616061.t0 vccd1.t15 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X152 a_350722_615130.t1 io_out[12].t0 a_350378_615130.t0 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=5.19 l=1.43
X153 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t11 a_343294_615747# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X154 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_345642_617070# vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X155 vccd1.t61 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t19 a_339370_613888.t13 vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X156 vccd1.t62 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t20 a_339370_613888.t12 vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X157 vccd1.t13 vccd1.t10 vccd1.t12 vccd1.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.258 ps=2.36 w=0.89 l=3.89
X158 a_335807_622237.t5 a_335719_622037.t9 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X159 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t3 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t14 a_341818_614929.t2 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X160 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t4 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_345642_614374.t5 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X161 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT a_345642_620402# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X162 gpio_analog[3].t4 a_341600_622217.t24 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X163 a_341818_619927.t0 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X164 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t13 a_345642_614374.t0 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X165 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t0 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg a_336716_619863# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X166 vccd1.t72 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t21 a_339370_617808# vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X167 vccd1.t1 a_336843_616061.t2 w_336471_617254# vccd1.t0 sky130_fd_pr__pfet_01v8 ad=0.687 pd=5.32 as=0.687 ps=5.32 w=2.37 l=4.38
X168 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_341818_618261.t0 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X169 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t3 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_345642_614374.t4 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X170 a_335719_622037.t1 a_335719_622037.t0 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X171 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t2 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_345642_614374.t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X172 vccd1.t73 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t22 a_339370_617808# vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X173 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT a_345642_621038.t6 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X174 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_345642_618736# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X175 a_345642_616040.t0 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X176 vccd1.t9 vccd1.t6 vccd1.t8 vccd1.t7 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=2
X177 a_341818_618261.t5 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t11 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X178 vccd1.t49 a_350378_615130.t4 io_out[15].t4 vccd1.t48 sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.9 as=1.5 ps=10.9 w=5.17 l=0.37
X179 a_336716_619863# pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=5
X180 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t12 a_341600_622217.t2 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
R8 vssa1 io_clamp_high[1] sky130_fd_pr__res_generic_m3 w=11 l=0.25
X181 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_345642_621038.t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X182 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_345642_616040.t4 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X183 gpio_analog[3].t3 a_341600_622217.t25 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X184 a_350722_615130.t2 io_out[12].t1 a_350378_615130.t1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=5.19 l=1.43
X185 a_337674_621712# a_335807_622237.t22 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t2 vccd1.t7 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X186 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t1 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t12 a_341818_616595.t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X187 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT vssa1 vssa1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X188 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t4 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_343294_620745# vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X189 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=1.48 ps=10.8 w=5.1 l=0.66
X190 a_350942_613328.t4 gpio_analog[7].t9 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X191 vccd1.t5 vccd1.t2 vccd1.t4 vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=2
X192 vccd1.t74 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t23 a_339370_613888.t11 vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X193 vccd1.t41 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t24 a_339370_618592# vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X194 vccd1.t42 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t25 a_339370_613888.t10 vccd1.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X195 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t0 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t14 a_343294_614081# vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X196 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_345642_616040.t3 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X197 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT a_345642_619372.t1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X198 a_345642_614374.t1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X199 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_345642_616040.t2 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X200 vccd1.t64 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t7 a_337674_621712# vccd1.t21 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X201 a_341600_622217.t9 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t13 vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X202 a_341818_616595.t0 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t13 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X203 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t0 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t14 a_341818_616595.t2 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X204 vccd1.t56 a_337443_613718.t4 a_337443_613718.t5 vccd1.t55 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
D0 io_out[11].t4 vccd1.t54 sky130_fd_pr__diode_pd2nw_05v5_lvt pj=2.6e+06 area=4.225e+11
X205 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t15 a_343294_614081# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X206 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_345642_619372.t0 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X207 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t14 a_341600_622217.t1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X208 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t12 a_343294_617413# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X209 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT vssa1 vssa1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X210 gpio_analog[3].t2 a_341600_622217.t26 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X211 vccd1.t45 a_350942_613328.t0 a_350942_613328.t1 vccd1.t44 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X212 a_350378_615130.t5 io_out[15].t3 sky130_fd_pr__cap_mim_m3_1 l=15 w=4
X213 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t15 a_343294_620745# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X214 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X215 w_336471_617254# w_336471_617254# vssa1 w_336471_617254# sky130_fd_pr__pfet_01v8_lvt ad=0.255 pd=2.34 as=0.255 ps=2.34 w=0.88 l=6.97
X216 vccd1.t58 a_352038_622652.t0 a_352038_622652.t1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.89
X217 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.725 ps=5.58 w=2.5 l=1
X218 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=1.48 ps=10.8 w=5.1 l=0.66
X219 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t13 a_341818_618261.t1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X220 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t16 a_341600_622217.t8 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X221 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_345642_620402# vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X222 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_345642_621038.t2 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X223 io_out[15].t1 io_out[16].t1 a_350722_615130.t3 io_out[15].t0 sky130_fd_pr__pfet_01v8_lvt ad=1.76 pd=12.7 as=1.76 ps=12.7 w=6.07 l=1.27
X224 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_345642_613738# vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X225 gpio_analog[3].t1 a_341600_622217.t27 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X226 vdda1 a_341600_622217.t28 gpio_analog[3].t16 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X227 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t17 a_341600_622217.t0 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X228 a_339370_613888.t0 a_335807_622237.t23 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t5 vccd1.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X229 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t14 a_343294_619079# vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X230 vssa1 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t15 a_341818_614929.t6 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X231 a_345642_619372.t5 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X232 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t15 a_343294_617413# vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
R9 vssa1 io_clamp_low[2] sky130_fd_pr__res_generic_m3 w=11 l=0.25
X233 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t0 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X234 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT vssa1 vssa1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X235 gpio_analog[3].t0 a_341600_622217.t29 vssa1 vssa1 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X236 a_343294_614081# pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t15 vdda1 vdda1 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
R10 a_337443_613718.n0 a_337443_613718.t4 37.8394
R11 a_337443_613718.n0 a_337443_613718.t2 37.8394
R12 a_337443_613718.t0 a_337443_613718.n0 12.0988
R13 a_337443_613718.n0 a_337443_613718.t3 11.4337
R14 a_337443_613718.n0 a_337443_613718.t1 11.428
R15 a_337443_613718.n0 a_337443_613718.t5 11.428
R16 vccd1.n93 vccd1.n61 23340
R17 vccd1.n93 vccd1.n62 23336.5
R18 vccd1.n144 vccd1.n61 23336.5
R19 vccd1.n144 vccd1.n62 23332.9
R20 vccd1.n126 vccd1.n64 9769.41
R21 vccd1.n126 vccd1.n65 9769.41
R22 vccd1.n142 vccd1.n65 9769.41
R23 vccd1.n142 vccd1.n64 9769.41
R24 vccd1.n25 vccd1.n23 7521.18
R25 vccd1.n34 vccd1.n25 7517.65
R26 vccd1.n35 vccd1.n23 7517.65
R27 vccd1.n35 vccd1.n34 7514.12
R28 vccd1.n56 vccd1.n50 5841.18
R29 vccd1.n56 vccd1.n51 5841.18
R30 vccd1.n58 vccd1.n50 5837.65
R31 vccd1.n58 vccd1.n51 5837.65
R32 vccd1.n152 vccd1.n150 5294.12
R33 vccd1.n152 vccd1.n46 5294.12
R34 vccd1.n156 vccd1.n46 3772.94
R35 vccd1.n150 vccd1.n44 3049.41
R36 vccd1.n19 vccd1.n18 2985.88
R37 vccd1.n16 vccd1.n14 2985.88
R38 vccd1.n160 vccd1.n44 1517.65
R39 vccd1.n14 vccd1.n13 949.587
R40 vccd1.n18 vccd1.n17 949.587
R41 vccd1.n128 vccd1.n127 843.169
R42 vccd1.n127 vccd1.n124 842.972
R43 vccd1.n160 vccd1.n159 727.059
R44 vccd1.n55 vccd1.n49 623.059
R45 vccd1.n59 vccd1.n49 622.683
R46 vccd1.n145 vccd1.n60 620.077
R47 vccd1.n154 vccd1.n153 564.707
R48 vccd1.n146 vccd1.n145 475.827
R49 vccd1.n55 vccd1.n54 467.954
R50 vccd1.n36 vccd1.n22 459.671
R51 vccd1.n37 vccd1.n36 452.519
R52 vccd1.n57 vccd1.t43 431.565
R53 vccd1.n153 vccd1.n149 406.414
R54 vccd1.t15 vccd1.n50 378.753
R55 vccd1.t67 vccd1.t32 367.363
R56 vccd1.t46 vccd1.t67 367.363
R57 vccd1.t65 vccd1.t44 367.363
R58 vccd1.t11 vccd1.t65 367.363
R59 vccd1.n155 vccd1.n154 344.031
R60 vccd1.n148 vccd1.n48 337.954
R61 vccd1.n2 vccd1.t54 330
R62 vccd1.n139 vccd1.n138 325.146
R63 vccd1.n102 vccd1.n101 323.012
R64 vccd1.n57 vccd1.t0 319.678
R65 vccd1.n15 vccd1.n11 318.495
R66 vccd1.n15 vccd1.n12 318.495
R67 vccd1.n86 vccd1.n85 314.729
R68 vccd1.t43 vccd1.n51 291.885
R69 vccd1.n20 vccd1.n12 282.247
R70 vccd1.n33 vccd1.n32 254.948
R71 vccd1.n140 vccd1.n139 251.107
R72 vccd1.n92 vccd1.n91 251.107
R73 vccd1.n67 vccd1.n66 250.353
R74 vccd1.n96 vccd1.n95 250.353
R75 vccd1.n101 vccd1.n100 248.095
R76 vccd1.n100 vccd1.n99 248.095
R77 vccd1.n99 vccd1.n98 248.095
R78 vccd1.n98 vccd1.n97 248.095
R79 vccd1.n97 vccd1.n96 248.095
R80 vccd1.n91 vccd1.n90 248.095
R81 vccd1.n90 vccd1.n89 248.095
R82 vccd1.n89 vccd1.n88 248.095
R83 vccd1.n88 vccd1.n87 248.095
R84 vccd1.n87 vccd1.n86 248.095
R85 vccd1.t32 vccd1.n23 232.912
R86 vccd1.n33 vccd1.n22 231.79
R87 vccd1.n34 vccd1.t11 213.075
R88 vccd1.n21 vccd1.n11 209.695
R89 vccd1.n152 vccd1.t50 202.427
R90 vccd1.t55 vccd1.n45 199.849
R91 vccd1.n151 vccd1.t55 195.214
R92 vccd1.t44 vccd1.n24 193.233
R93 vccd1.t50 vccd1.n151 192.995
R94 vccd1.n148 vccd1.n59 189.365
R95 vccd1.n26 vccd1.n9 186.632
R96 vccd1.n24 vccd1.t46 174.131
R97 vccd1.n66 vccd1.n60 162.636
R98 vccd1.n112 vccd1.n108 150.589
R99 vccd1.n106 vccd1.n102 150.589
R100 vccd1.n85 vccd1.n81 150.589
R101 vccd1.n79 vccd1.n75 150.589
R102 vccd1.t25 vccd1.n143 141.708
R103 vccd1.n54 vccd1.n53 138.542
R104 vccd1.n75 vccd1.n74 133.732
R105 vccd1.n94 vccd1.n92 127.624
R106 vccd1.n141 vccd1.n140 126.118
R107 vccd1.n141 vccd1.n67 121.977
R108 vccd1.n95 vccd1.n94 120.472
R109 vccd1.n126 vccd1.t7 119.335
R110 vccd1.n116 vccd1.n71 107.016
R111 vccd1.n116 vccd1.n115 107.016
R112 vccd1.n122 vccd1.n70 107.016
R113 vccd1.n122 vccd1.n121 107.016
R114 vccd1.n130 vccd1.n69 107.016
R115 vccd1.n130 vccd1.n129 107.016
R116 vccd1.n136 vccd1.n68 107.016
R117 vccd1.n136 vccd1.n135 107.016
R118 vccd1.n125 vccd1.t21 96.026
R119 vccd1.n111 vccd1.t27 94.1656
R120 vccd1.n109 vccd1.t26 94.1656
R121 vccd1.n105 vccd1.t5 94.1656
R122 vccd1.n103 vccd1.t4 94.1656
R123 vccd1.n84 vccd1.t29 94.1656
R124 vccd1.n82 vccd1.t30 94.1656
R125 vccd1.n78 vccd1.t39 94.1656
R126 vccd1.n76 vccd1.t40 94.1656
R127 vccd1.n143 vccd1.t21 90.4323
R128 vccd1.n73 vccd1.n72 82.4476
R129 pmu_circuits_0.iref_2nA_0.iref_2nA_vref_0.DD vccd1.n147 80.1379
R130 vccd1.n39 vccd1.n10 75.614
R131 vccd1.n110 vccd1.n109 75.2946
R132 vccd1.n111 vccd1.n110 75.2946
R133 vccd1.n104 vccd1.n103 75.2946
R134 vccd1.n105 vccd1.n104 75.2946
R135 vccd1.n84 vccd1.n83 75.2946
R136 vccd1.n83 vccd1.n82 75.2946
R137 vccd1.n78 vccd1.n77 75.2946
R138 vccd1.n77 vccd1.n76 75.2946
R139 vccd1.t7 vccd1.n125 67.1251
R140 vccd1.n134 vccd1.n133 64.6279
R141 vccd1.n119 vccd1.n118 64.4315
R142 vccd1.n38 vccd1.n21 63.0245
R143 vccd1.n114 vccd1.n113 62.5491
R144 vccd1.n22 vccd1.t13 60.0995
R145 vccd1.n37 vccd1.t34 60.0995
R146 vccd1.n144 vccd1.t25 59.4732
R147 vccd1.n113 vccd1.n112 58.6643
R148 vccd1.n93 vccd1.t3 58.3834
R149 vccd1.n115 vccd1.t36 57.1406
R150 vccd1.n71 vccd1.t37 57.1406
R151 vccd1.n121 vccd1.t18 57.1406
R152 vccd1.n70 vccd1.t19 57.1406
R153 vccd1.n129 vccd1.t9 57.1406
R154 vccd1.n69 vccd1.t8 57.1406
R155 vccd1.n135 vccd1.t23 57.1406
R156 vccd1.n68 vccd1.t22 57.1406
R157 vccd1.n52 vccd1.t16 57.1406
R158 vccd1.n38 vccd1.n37 53.4946
R159 vccd1.n32 vccd1.t12 48.3828
R160 vccd1.n26 vccd1.t33 45.276
R161 vccd1.n53 vccd1.n48 45.1973
R162 vccd1.n107 vccd1.n106 40.6593
R163 vccd1.n81 vccd1.n80 40.6593
R164 vccd1.n108 vccd1.n107 37.6476
R165 vccd1.n80 vccd1.n79 37.6476
R166 vccd1.n28 vccd1.n27 34.174
R167 vccd1.n31 vccd1.n30 34.174
R168 vccd1.n54 vccd1.n52 33.746
R169 vccd1.n112 vccd1.n111 32.8353
R170 vccd1.n109 vccd1.n108 32.8353
R171 vccd1.n106 vccd1.n105 32.8353
R172 vccd1.n103 vccd1.n102 32.8353
R173 vccd1.n31 vccd1.t66 32.0995
R174 vccd1.n30 vccd1.t45 32.0995
R175 vccd1.n28 vccd1.t47 32.0995
R176 vccd1.n27 vccd1.t68 32.0995
R177 vccd1.n27 vccd1.n26 28.5054
R178 vccd1.n32 vccd1.n31 28.5054
R179 vccd1.t3 vccd1.n63 28.2824
R180 vccd1.n139 vccd1.t63 27.7091
R181 vccd1.n140 vccd1.t76 27.7091
R182 vccd1.n67 vccd1.t75 27.7091
R183 vccd1.n66 vccd1.t64 27.7091
R184 vccd1.t25 vccd1.n63 27.6433
R185 vccd1.n118 vccd1.n71 26.9918
R186 vccd1.n115 vccd1.n114 26.9918
R187 vccd1.n124 vccd1.n70 26.9918
R188 vccd1.n121 vccd1.n120 26.9918
R189 vccd1.n132 vccd1.n69 26.9918
R190 vccd1.n129 vccd1.n128 26.9918
R191 vccd1.n138 vccd1.n68 26.9918
R192 vccd1.n135 vccd1.n134 26.9918
R193 vccd1.n85 vccd1.n84 26.4353
R194 vccd1.n82 vccd1.n81 26.4353
R195 vccd1.n79 vccd1.n78 26.4353
R196 vccd1.n76 vccd1.n75 26.4353
R197 vccd1.n101 vccd1.t51 26.3779
R198 vccd1.n100 vccd1.t60 26.3779
R199 vccd1.n99 vccd1.t61 26.3779
R200 vccd1.n98 vccd1.t74 26.3779
R201 vccd1.n97 vccd1.t70 26.3779
R202 vccd1.n96 vccd1.t73 26.3779
R203 vccd1.n95 vccd1.t52 26.3779
R204 vccd1.n92 vccd1.t41 26.3779
R205 vccd1.n91 vccd1.t72 26.3779
R206 vccd1.n90 vccd1.t69 26.3779
R207 vccd1.n89 vccd1.t62 26.3779
R208 vccd1.n88 vccd1.t42 26.3779
R209 vccd1.n87 vccd1.t71 26.3779
R210 vccd1.n86 vccd1.t53 26.3779
R211 vccd1.t0 vccd1.t15 25.0188
R212 vccd1.n74 vccd1.n47 21.3338
R213 vccd1.n132 vccd1.n131 20.6846
R214 vccd1.n131 vccd1.n128 20.6846
R215 vccd1.n138 vccd1.n137 20.6846
R216 vccd1.n137 vccd1.n134 20.6846
R217 vccd1.n117 vccd1.n114 18.7794
R218 vccd1.n118 vccd1.n117 18.7794
R219 vccd1.n123 vccd1.n120 18.7794
R220 vccd1.n124 vccd1.n123 18.7794
R221 vccd1.n30 vccd1.n29 18.0327
R222 vccd1.n133 vccd1.n132 17.9456
R223 vccd1.n120 vccd1.n119 17.7491
R224 vccd1.n42 vccd1.t56 17.5661
R225 vccd1.n147 vccd1.n146 17.4227
R226 vccd1.n29 vccd1.n28 16.1418
R227 vccd1.n77 vccd1.t38 13.7387
R228 vccd1.n83 vccd1.t28 13.7387
R229 vccd1.n104 vccd1.t2 13.7387
R230 vccd1.n110 vccd1.t24 13.7387
R231 vccd1.n117 vccd1.t35 13.7387
R232 vccd1.t35 vccd1.n116 13.7387
R233 vccd1.n123 vccd1.t17 13.7387
R234 vccd1.t17 vccd1.n122 13.7387
R235 vccd1.n131 vccd1.t6 13.7387
R236 vccd1.t6 vccd1.n130 13.7387
R237 vccd1.n137 vccd1.t20 13.7387
R238 vccd1.t20 vccd1.n136 13.7387
R239 vccd1.n113 vccd1.n60 13.6867
R240 vccd1.n160 vccd1.n45 13.4821
R241 vccd1.n72 vccd1.n47 13.177
R242 vccd1.n48 vccd1.t1 12.0543
R243 vccd1.n72 vccd1.t57 11.4275
R244 vccd1.n21 vccd1.n20 10.8113
R245 pmu_circuits_0.iref_2nA_0.DD vccd1.n161 10.2882
R246 vccd1.n10 vccd1.t31 9.47999
R247 vccd1.n33 vccd1.t10 9.47999
R248 vccd1.n7 vccd1.n6 9.3005
R249 vccd1.n161 vccd1.n160 8.85536
R250 vccd1.n148 pmu_circuits_0.iref_2nA_0.iref_2nA_vref_0.DD 8.72328
R251 vccd1.n39 vccd1.n38 8.40959
R252 vccd1.n40 vccd1.n9 8.10924
R253 vccd1.n20 vccd1.t49 5.52608
R254 vccd1.n40 vccd1.n39 5.40633
R255 pmu_circuits_0.vref01_0.DD vccd1.t59 4.9842
R256 vccd1.n146 vccd1.n42 4.44294
R257 vccd1.n1 vccd1.t58 4.3481
R258 vccd1.n161 vccd1.n43 4.28102
R259 vccd1.n52 vccd1.t14 4.11799
R260 vccd1.n161 vccd1.n42 3.88459
R261 pmu_circuits_0.dd_01 vccd1.n0 3.61179
R262 vccd1.n3 vccd1.n2 2.84494
R263 vccd1 vccd1.n43 2.82647
R264 vccd1.n5 vccd1.n4 2.8192
R265 vccd1.n162 pmu_circuits_0.iref_2nA_0.DD 2.56417
R266 vccd1.n149 vccd1.n148 2.44683
R267 vccd1.n162 vccd1.n41 2.08208
R268 vccd1.n41 pmu_circuits_0.ldo_0.DD 1.29471
R269 vccd1.n41 vccd1.n8 1.26929
R270 vccd1.n8 vccd1.n7 1.17606
R271 vccd1.n8 vccd1.n1 1.01403
R272 vccd1.n155 vccd1.n47 0.970197
R273 vccd1.n10 vccd1.n9 0.840904
R274 pmu_circuits_0.dd_01 vccd1.n162 0.758737
R275 vccd1.n74 vccd1.n73 0.706994
R276 vccd1.n73 vccd1 0.644656
R277 vccd1.n157 vccd1.n45 0.28389
R278 pmu_circuits_0.ldo_0.DD vccd1.n40 0.196382
R279 vccd1.n0 vccd1 0.183467
R280 vccd1.n0 VCCD1 0.155422
R281 vccd1.n7 vccd1.n5 0.115443
R282 VCCD1 vccd1 0.100257
R283 vccd1.n1 pmu_circuits_0.vref01_0.DD 0.0587192
R284 vccd1.n147 vccd1.n44 0.0402849
R285 vccd1.n157 vccd1.n44 0.0402849
R286 vccd1.n14 vccd1.n11 0.025954
R287 vccd1.n18 vccd1.n12 0.025954
R288 vccd1.n158 vccd1.n156 0.0146429
R289 vccd1.n156 vccd1.n155 0.0141431
R290 vccd1.n159 vccd1.n158 0.00674884
R291 vccd1.n159 vccd1.n43 0.00624891
R292 vccd1.n34 vccd1.n33 0.00450849
R293 vccd1.n23 vccd1.n10 0.00450849
R294 vccd1.n51 vccd1.n49 0.00424858
R295 vccd1.n53 vccd1.n50 0.00424858
R296 vccd1.n16 vccd1.n15 0.00414317
R297 vccd1.n20 vccd1.n19 0.00414317
R298 vccd1.n150 vccd1.n149 0.00377503
R299 vccd1.n151 vccd1.n150 0.00377503
R300 vccd1.n154 vccd1.n46 0.00377503
R301 vccd1.n151 vccd1.n46 0.00377503
R302 vccd1.n107 vccd1.n61 0.00369903
R303 vccd1.n63 vccd1.n61 0.00369903
R304 vccd1.n63 vccd1.n62 0.00369903
R305 vccd1.n80 vccd1.n62 0.00369903
R306 vccd1.n19 vccd1.n13 0.00355895
R307 vccd1.n17 vccd1.n16 0.00348454
R308 vccd1.n119 vccd1.n64 0.00338999
R309 vccd1.n125 vccd1.n64 0.00338999
R310 vccd1.n125 vccd1.n65 0.00338999
R311 vccd1.n133 vccd1.n65 0.00338999
R312 vccd1.n153 vccd1.n152 0.00337446
R313 vccd1.n56 vccd1.n55 0.00268001
R314 vccd1.n57 vccd1.n56 0.00268001
R315 vccd1.n59 vccd1.n58 0.00268001
R316 vccd1.n58 vccd1.n57 0.00268001
R317 vccd1.t48 vccd1.n13 0.00231816
R318 vccd1.n17 vccd1.t48 0.00215862
R319 vccd1.n29 vccd1.n25 0.00193193
R320 vccd1.n25 vccd1.n24 0.00193193
R321 vccd1.n35 vccd1.n24 0.00193193
R322 vccd1.n36 vccd1.n35 0.00193193
R323 vccd1.n127 vccd1.n126 0.00161095
R324 vccd1.n142 vccd1.n141 0.00161095
R325 vccd1.n143 vccd1.n142 0.00161095
R326 vccd1.n158 vccd1.n157 0.00100005
R327 vccd1.n145 vccd1.n144 0.000866167
R328 vccd1.n94 vccd1.n93 0.000866167
R329 vccd1.n5 vccd1.n3 0.00051539
R330 a_335807_622237.t9 a_335807_622237.n2 151.024
R331 a_335807_622237.t21 a_335807_622237.t15 75.728
R332 a_335807_622237.t12 a_335807_622237.t9 75.728
R333 a_335807_622237.t13 a_335807_622237.t12 75.728
R334 a_335807_622237.t18 a_335807_622237.t13 75.728
R335 a_335807_622237.t6 a_335807_622237.t18 75.728
R336 a_335807_622237.t17 a_335807_622237.t6 75.728
R337 a_335807_622237.t10 a_335807_622237.t17 75.728
R338 a_335807_622237.t19 a_335807_622237.t10 75.728
R339 a_335807_622237.t16 a_335807_622237.t19 75.728
R340 a_335807_622237.t23 a_335807_622237.t16 75.728
R341 a_335807_622237.t14 a_335807_622237.t23 75.728
R342 a_335807_622237.t20 a_335807_622237.t14 75.728
R343 a_335807_622237.t8 a_335807_622237.t20 75.728
R344 a_335807_622237.t11 a_335807_622237.t8 75.728
R345 a_335807_622237.t15 a_335807_622237.t7 73.0385
R346 a_335807_622237.n2 a_335807_622237.t21 61.9359
R347 a_335807_622237.n1 a_335807_622237.t11 41.3671
R348 a_335807_622237.n0 a_335807_622237.t2 37.8394
R349 a_335807_622237.n0 a_335807_622237.t0 37.8394
R350 a_335807_622237.n3 a_335807_622237.t5 13.5808
R351 a_335807_622237.n4 a_335807_622237.t1 11.428
R352 a_335807_622237.t3 a_335807_622237.n5 11.428
R353 a_335807_622237.n2 a_335807_622237.t22 11.0702
R354 a_335807_622237.n3 a_335807_622237.t4 10.6813
R355 a_335807_622237.n1 a_335807_622237.n3 7.30437
R356 a_335807_622237.n4 a_335807_622237.n1 0.573403
R357 a_335807_622237.n0 a_335807_622237.n4 0.555619
R358 a_335807_622237.n5 a_335807_622237.n0 0.403391
R359 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t18 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t15 75.728
R360 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t19 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t18 75.728
R361 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t23 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t19 75.728
R362 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t13 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t23 75.728
R363 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t22 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t13 75.728
R364 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t16 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t22 75.728
R365 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t24 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t16 75.728
R366 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t21 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t24 75.728
R367 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t12 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t21 75.728
R368 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t20 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t12 75.728
R369 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t25 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t20 75.728
R370 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t14 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t25 75.728
R371 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n6 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t17 37.8646
R372 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n6 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t14 37.8639
R373 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n4 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t5 12.8247
R374 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n5 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t2 12.8247
R375 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n2 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t3 12.8247
R376 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n3 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t8 12.8247
R377 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n0 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t6 11.428
R378 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n4 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t9 11.428
R379 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n5 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t4 11.428
R380 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t10 11.428
R381 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n2 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t11 11.428
R382 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n3 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t7 11.428
R383 pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Ip2 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n1 8.50055
R384 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n7 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t0 8.17163
R385 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t1 7.50959
R386 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n7 pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Ip2 5.32175
R387 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n7 3.49672
R388 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n0 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n6 2.74398
R389 pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Ip2 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n0 0.990509
R390 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n0 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n5 0.810482
R391 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n3 0.810433
R392 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n0 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n4 0.810432
R393 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n2 0.810432
R394 a_339370_613888.n1 a_339370_613888.t18 11.554
R395 a_339370_613888.n0 a_339370_613888.t19 11.554
R396 a_339370_613888.n6 a_339370_613888.t15 11.554
R397 a_339370_613888.n7 a_339370_613888.t17 11.554
R398 a_339370_613888.n8 a_339370_613888.t10 11.554
R399 a_339370_613888.n9 a_339370_613888.t12 11.554
R400 a_339370_613888.n2 a_339370_613888.t16 11.554
R401 a_339370_613888.n3 a_339370_613888.t14 11.554
R402 a_339370_613888.n4 a_339370_613888.t13 11.554
R403 a_339370_613888.n5 a_339370_613888.t11 11.554
R404 a_339370_613888.n0 a_339370_613888.t0 11.5402
R405 a_339370_613888.n6 a_339370_613888.t6 11.5402
R406 a_339370_613888.n7 a_339370_613888.t8 11.5402
R407 a_339370_613888.n8 a_339370_613888.t1 11.5402
R408 a_339370_613888.n9 a_339370_613888.t3 11.5402
R409 a_339370_613888.n2 a_339370_613888.t7 11.5402
R410 a_339370_613888.n3 a_339370_613888.t5 11.5402
R411 a_339370_613888.n4 a_339370_613888.t4 11.5402
R412 a_339370_613888.n5 a_339370_613888.t2 11.5402
R413 a_339370_613888.t9 a_339370_613888.n1 11.5402
R414 a_339370_613888.n1 a_339370_613888.n0 7.86782
R415 a_339370_613888.n7 a_339370_613888.n6 1.26396
R416 a_339370_613888.n8 a_339370_613888.n7 1.26396
R417 a_339370_613888.n9 a_339370_613888.n8 1.26396
R418 a_339370_613888.n3 a_339370_613888.n2 1.26396
R419 a_339370_613888.n4 a_339370_613888.n3 1.26396
R420 a_339370_613888.n5 a_339370_613888.n4 1.26396
R421 a_339370_613888.n1 a_339370_613888.n5 1.26396
R422 a_339370_613888.n0 a_339370_613888.n9 1.26396
R423 a_350942_613328.n0 a_350942_613328.t1 32.4466
R424 a_350942_613328.n0 a_350942_613328.t3 32.4466
R425 a_350942_613328.t0 a_350942_613328.t6 19.1411
R426 a_350942_613328.t2 a_350942_613328.t7 19.1411
R427 a_350942_613328.n3 a_350942_613328.t5 10.1828
R428 a_350942_613328.n2 a_350942_613328.t0 9.48031
R429 a_350942_613328.n1 a_350942_613328.t2 9.48031
R430 a_350942_613328.n3 a_350942_613328.n0 5.92365
R431 a_350942_613328.t4 a_350942_613328.n3 5.36911
R432 a_350942_613328.n0 a_350942_613328.n2 0.450838
R433 a_350942_613328.n0 a_350942_613328.n1 0.351043
R434 a_350378_615130.n0 a_350378_615130.t4 191.636
R435 a_350378_615130.n0 a_350378_615130.t3 34.661
R436 a_350378_615130.n0 a_350378_615130.t2 33.291
R437 a_350378_615130.n2 a_350378_615130.t1 4.51459
R438 a_350378_615130.t0 a_350378_615130.n2 3.35375
R439 a_350378_615130.n1 a_350378_615130.n0 2.51069
R440 a_350378_615130.n2 a_350378_615130.n1 1.37236
R441 a_350378_615130.n1 a_350378_615130.t5 0.251842
R442 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n0 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t6 21.4396
R443 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n0 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t5 18.8004
R444 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t4 18.8004
R445 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n2 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t7 18.8004
R446 pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Ip1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t3 11.5886
R447 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n3 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t2 11.5885
R448 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n4 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t0 8.4133
R449 pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Ip1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n2 7.65117
R450 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t1 7.50959
R451 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n3 pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Ip1 3.82182
R452 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n0 2.63976
R453 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n2 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n1 2.63976
R454 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n4 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n3 1.93205
R455 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n4 0.573
R456 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n17 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t4 265.382
R457 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n19 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n18 262.217
R458 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n7 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t12 183.099
R459 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n6 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t6 183.099
R460 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t6 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n5 183.099
R461 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n2 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t8 182.653
R462 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t12 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n0 182.297
R463 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n2 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t11 182.288
R464 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n1 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t14 182.285
R465 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n6 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t7 182.263
R466 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t14 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n7 182.263
R467 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t7 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n5 182.263
R468 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n18 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t1 155.667
R469 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n17 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t0 155.667
R470 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t9 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n4 146.282
R471 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t13 145.889
R472 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t13 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n10 145.857
R473 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n8 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t9 145.851
R474 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n12 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t5 135.911
R475 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n15 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n14 122.928
R476 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n18 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n17 109.715
R477 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t15 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n13 98.2234
R478 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n15 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t15 49.4098
R479 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n3 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t10 45.8204
R480 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n12 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n3 28.5785
R481 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n14 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t2 28.5685
R482 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t5 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n11 19.7637
R483 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n16 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n15 5.00095
R484 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n9 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n4 4.13208
R485 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n19 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t3 3.16453
R486 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n16 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n2 1.3453
R487 pmu_circuits_0.ring_100mV_0.mdls_inv_8.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n19 1.29092
R488 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n13 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n12 1.06388
R489 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n7 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n6 0.835457
R490 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n1 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n5 0.813812
R491 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n1 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n0 0.810242
R492 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n10 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n9 0.607643
R493 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n4 0.454134
R494 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n9 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n8 0.43198
R495 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n11 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN 0.339159
R496 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n8 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n1 0.320167
R497 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n10 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n0 0.21421
R498 pmu_circuits_0.ring_100mV_0.mdls_inv_8.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n16 0.184521
R499 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n17 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n9 368.413
R500 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n22 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t0 265.382
R501 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n24 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n23 262.217
R502 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n10 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t10 251.451
R503 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t15 182.653
R504 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t8 182.288
R505 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n10 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t17 182.262
R506 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n11 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t14 182.262
R507 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n12 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t12 182.262
R508 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n13 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t6 182.262
R509 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n14 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t5 182.262
R510 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n15 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t9 182.262
R511 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n16 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t7 182.262
R512 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n23 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t3 155.667
R513 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n22 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t2 155.667
R514 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n20 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n19 122.928
R515 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n23 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n22 109.715
R516 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t11 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n18 98.2234
R517 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n9 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n8 72.1132
R518 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n8 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n7 72.1132
R519 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n7 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n6 72.1132
R520 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n6 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n5 72.1132
R521 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n5 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n4 72.1132
R522 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n4 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n3 72.1132
R523 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n16 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n15 69.1897
R524 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n15 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n14 69.1897
R525 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n14 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n13 69.1897
R526 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n13 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n12 69.1897
R527 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n12 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n11 69.1897
R528 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n11 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n10 69.1897
R529 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n17 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n16 62.0129
R530 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n20 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t11 49.4098
R531 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n2 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t13 36.7438
R532 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n2 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t16 32.5647
R533 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n19 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t4 28.5685
R534 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n0 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n17 27.9962
R535 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n0 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n2 6.45024
R536 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n21 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n20 5.00095
R537 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n24 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t1 3.16453
R538 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n18 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n0 2.08823
R539 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n21 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n1 1.3453
R540 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n24 1.29092
R541 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n21 0.184521
R542 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n0 pmu_circuits_0.ring_100mV_0.ring_100mV_buffer_0.IN 0.156641
R543 a_341600_622217.n25 a_341600_622217.t14 332.849
R544 a_341600_622217.n5 a_341600_622217.n4 212.389
R545 a_341600_622217.n5 a_341600_622217.t19 182.262
R546 a_341600_622217.n6 a_341600_622217.t16 182.262
R547 a_341600_622217.n7 a_341600_622217.t13 182.262
R548 a_341600_622217.n8 a_341600_622217.t21 182.262
R549 a_341600_622217.n9 a_341600_622217.t20 182.262
R550 a_341600_622217.n16 a_341600_622217.t24 182.262
R551 a_341600_622217.t24 a_341600_622217.n15 182.262
R552 a_341600_622217.n17 a_341600_622217.t23 182.262
R553 a_341600_622217.n20 a_341600_622217.t22 182.262
R554 a_341600_622217.t22 a_341600_622217.n19 182.262
R555 a_341600_622217.n21 a_341600_622217.t26 182.262
R556 a_341600_622217.n24 a_341600_622217.t25 182.262
R557 a_341600_622217.t25 a_341600_622217.n23 182.262
R558 a_341600_622217.n32 a_341600_622217.t12 182.262
R559 a_341600_622217.t12 a_341600_622217.n31 182.262
R560 a_341600_622217.n27 a_341600_622217.t10 182.262
R561 a_341600_622217.n26 a_341600_622217.t27 182.262
R562 a_341600_622217.n25 a_341600_622217.t17 182.262
R563 a_341600_622217.n29 a_341600_622217.n28 150.589
R564 a_341600_622217.n30 a_341600_622217.n29 150.589
R565 a_341600_622217.n31 a_341600_622217.n30 150.589
R566 a_341600_622217.n23 a_341600_622217.n22 150.589
R567 a_341600_622217.n19 a_341600_622217.n18 150.589
R568 a_341600_622217.n15 a_341600_622217.n14 150.589
R569 a_341600_622217.n14 a_341600_622217.n13 150.589
R570 a_341600_622217.n13 a_341600_622217.n12 150.589
R571 a_341600_622217.n12 a_341600_622217.n11 150.589
R572 a_341600_622217.n11 a_341600_622217.n10 150.589
R573 a_341600_622217.n24 a_341600_622217.n21 150.589
R574 a_341600_622217.n21 a_341600_622217.n20 150.589
R575 a_341600_622217.n20 a_341600_622217.n17 150.589
R576 a_341600_622217.n17 a_341600_622217.n16 150.589
R577 a_341600_622217.n16 a_341600_622217.n9 150.589
R578 a_341600_622217.n9 a_341600_622217.n8 150.589
R579 a_341600_622217.n8 a_341600_622217.n7 150.589
R580 a_341600_622217.n7 a_341600_622217.n6 150.589
R581 a_341600_622217.n6 a_341600_622217.n5 150.589
R582 a_341600_622217.n26 a_341600_622217.n25 150.589
R583 a_341600_622217.n27 a_341600_622217.n26 150.589
R584 a_341600_622217.n32 a_341600_622217.n27 150.589
R585 a_341600_622217.n36 a_341600_622217.n35 150.589
R586 a_341600_622217.n38 a_341600_622217.n37 150.589
R587 a_341600_622217.n35 a_341600_622217.n34 96.6009
R588 a_341600_622217.n40 a_341600_622217.n39 87.4672
R589 a_341600_622217.n40 a_341600_622217.n36 66.2593
R590 a_341600_622217.n39 a_341600_622217.n38 66.2593
R591 a_341600_622217.n41 a_341600_622217.n40 66.2593
R592 a_341600_622217.n36 a_341600_622217.t28 49.4098
R593 a_341600_622217.n35 a_341600_622217.t18 49.4098
R594 a_341600_622217.n41 a_341600_622217.t11 49.4098
R595 a_341600_622217.n33 a_341600_622217.n32 46.6829
R596 a_341600_622217.n34 a_341600_622217.t15 42.6645
R597 a_341600_622217.n4 a_341600_622217.t29 40.6427
R598 a_341600_622217.n33 a_341600_622217.n24 38.777
R599 a_341600_622217.n43 a_341600_622217.n33 32.5457
R600 a_341600_622217.n43 a_341600_622217.t8 30.2238
R601 a_341600_622217.n42 a_341600_622217.t9 28.5701
R602 a_341600_622217.n0 a_341600_622217.t3 5.95384
R603 a_341600_622217.n44 a_341600_622217.n43 4.84496
R604 a_341600_622217.n44 a_341600_622217.t5 4.60076
R605 a_341600_622217.n45 a_341600_622217.t4 4.60076
R606 a_341600_622217.n0 a_341600_622217.t0 4.59778
R607 a_341600_622217.n1 a_341600_622217.t1 4.59778
R608 a_341600_622217.n2 a_341600_622217.t2 4.59778
R609 a_341600_622217.n3 a_341600_622217.t6 4.59778
R610 a_341600_622217.t7 a_341600_622217.n46 4.59778
R611 a_341600_622217.n43 a_341600_622217.n42 2.10396
R612 a_341600_622217.n42 a_341600_622217.n41 1.96379
R613 a_341600_622217.n1 a_341600_622217.n0 1.35656
R614 a_341600_622217.n2 a_341600_622217.n1 1.35656
R615 a_341600_622217.n3 a_341600_622217.n2 1.35656
R616 a_341600_622217.n46 a_341600_622217.n3 1.35656
R617 a_341600_622217.n46 a_341600_622217.n45 1.33027
R618 a_341600_622217.n45 a_341600_622217.n44 1.31668
R619 gpio_analog[3].n19 gpio_analog[3] 222.178
R620 gpio_analog[3].n0 gpio_analog[3].t19 30.4433
R621 gpio_analog[3].n2 gpio_analog[3].t18 29.7591
R622 gpio_analog[3].n0 gpio_analog[3].t16 29.2657
R623 gpio_analog[3].n1 gpio_analog[3].t17 29.2657
R624 gpio_analog[3].n4 gpio_analog[3].t0 5.86456
R625 gpio_analog[3] gpio_analog[3].t12 4.50884
R626 gpio_analog[3].n4 gpio_analog[3].t9 4.5085
R627 gpio_analog[3].n5 gpio_analog[3].t11 4.5085
R628 gpio_analog[3].n6 gpio_analog[3].t13 4.5085
R629 gpio_analog[3].n7 gpio_analog[3].t7 4.5085
R630 gpio_analog[3].n8 gpio_analog[3].t8 4.5085
R631 gpio_analog[3].n9 gpio_analog[3].t4 4.5085
R632 gpio_analog[3].n10 gpio_analog[3].t5 4.5085
R633 gpio_analog[3].n11 gpio_analog[3].t6 4.5085
R634 gpio_analog[3].n12 gpio_analog[3].t2 4.5085
R635 gpio_analog[3].n13 gpio_analog[3].t3 4.5085
R636 gpio_analog[3].n14 gpio_analog[3].t14 4.5085
R637 gpio_analog[3].n15 gpio_analog[3].t15 4.5085
R638 gpio_analog[3].n17 gpio_analog[3].t10 4.4579
R639 gpio_analog[3].n16 gpio_analog[3].t1 4.4579
R640 gpio_analog[3].n1 gpio_analog[3].n0 2.18471
R641 gpio_analog[3].n19 gpio_analog[3].n18 1.87736
R642 gpio_analog[3].n5 gpio_analog[3].n4 1.35656
R643 gpio_analog[3].n6 gpio_analog[3].n5 1.35656
R644 gpio_analog[3].n7 gpio_analog[3].n6 1.35656
R645 gpio_analog[3].n8 gpio_analog[3].n7 1.35656
R646 gpio_analog[3].n9 gpio_analog[3].n8 1.35656
R647 gpio_analog[3].n10 gpio_analog[3].n9 1.35656
R648 gpio_analog[3].n11 gpio_analog[3].n10 1.35656
R649 gpio_analog[3].n12 gpio_analog[3].n11 1.35656
R650 gpio_analog[3].n13 gpio_analog[3].n12 1.35656
R651 gpio_analog[3].n14 gpio_analog[3].n13 1.35656
R652 gpio_analog[3].n15 gpio_analog[3].n14 1.35656
R653 gpio_analog[3].n16 gpio_analog[3].n15 0.685584
R654 gpio_analog[3].n2 gpio_analog[3].n1 0.303132
R655 gpio_analog[3].n3 gpio_analog[3].n2 0.221405
R656 gpio_analog[3].n17 gpio_analog[3].n16 0.15724
R657 gpio_analog[3].n19 pmu_circuits_0.ring_out 0.102583
R658 gpio_analog[3].n18 gpio_analog[3].n3 0.0490893
R659 gpio_analog[3].n3 gpio_analog[3] 0.0463464
R660 pmu_circuits_0.ring_out gpio_analog[3].n19 0.0284412
R661 gpio_analog[3].n18 gpio_analog[3].n17 0.0118636
R662 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n17 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t4 265.382
R663 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n19 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n18 262.217
R664 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n7 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t7 183.099
R665 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n6 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t14 183.099
R666 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t14 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n5 183.099
R667 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n2 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t15 182.653
R668 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t7 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n0 182.297
R669 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n2 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t6 182.288
R670 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n1 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t11 182.285
R671 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n6 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t9 182.263
R672 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t11 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n7 182.263
R673 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t9 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n5 182.263
R674 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n17 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t2 155.667
R675 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n18 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t1 155.667
R676 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t5 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n4 146.282
R677 pmu_circuits_0.ring_100mV_0.mdls_inv_8.IN pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t10 145.889
R678 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t10 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n10 145.857
R679 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n8 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t5 145.851
R680 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n12 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t8 135.911
R681 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n15 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n14 122.928
R682 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n18 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n17 109.715
R683 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t13 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n13 98.2234
R684 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n15 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t13 49.4098
R685 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n3 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t12 45.8204
R686 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n12 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n3 28.5785
R687 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n14 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t0 28.5685
R688 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t8 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n11 19.7637
R689 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n16 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n15 5.00095
R690 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n9 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n4 4.13208
R691 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n19 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t3 3.16453
R692 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n13 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n12 2.84116
R693 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n16 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n2 1.3453
R694 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n19 1.29092
R695 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n7 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n6 0.835457
R696 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n1 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n5 0.813812
R697 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n1 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n0 0.810242
R698 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n10 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n9 0.607643
R699 pmu_circuits_0.ring_100mV_0.mdls_inv_8.IN pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n4 0.454134
R700 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n9 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n8 0.43198
R701 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n11 pmu_circuits_0.ring_100mV_0.mdls_inv_8.IN 0.339159
R702 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n8 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n1 0.320167
R703 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n10 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n0 0.21421
R704 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n16 0.184521
R705 a_341818_614929.n1 a_341818_614929.t2 260.2
R706 a_341818_614929.n0 a_341818_614929.t6 252.136
R707 a_341818_614929.t5 a_341818_614929.n4 251.333
R708 a_341818_614929.n2 a_341818_614929.n0 164.748
R709 a_341818_614929.n4 a_341818_614929.t0 157.893
R710 a_341818_614929.n3 a_341818_614929.t3 155.667
R711 a_341818_614929.n1 a_341818_614929.t4 149.827
R712 a_341818_614929.n3 a_341818_614929.n2 72.9605
R713 a_341818_614929.n2 a_341818_614929.n1 9.14336
R714 a_341818_614929.n4 a_341818_614929.n3 8.74717
R715 a_341818_614929.n0 a_341818_614929.t1 3.16453
R716 a_341818_616595.n2 a_341818_616595.t5 260.2
R717 a_341818_616595.n4 a_341818_616595.t6 252.136
R718 a_341818_616595.n0 a_341818_616595.t3 251.333
R719 a_341818_616595.n4 a_341818_616595.n3 164.748
R720 a_341818_616595.n0 a_341818_616595.t0 157.893
R721 a_341818_616595.n1 a_341818_616595.t2 155.667
R722 a_341818_616595.n2 a_341818_616595.t4 149.827
R723 a_341818_616595.n3 a_341818_616595.n1 72.9605
R724 a_341818_616595.n3 a_341818_616595.n2 9.14336
R725 a_341818_616595.n1 a_341818_616595.n0 8.74717
R726 a_341818_616595.t1 a_341818_616595.n4 3.16453
R727 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n19 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t1 265.382
R728 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n21 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n20 262.217
R729 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n6 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t13 183.099
R730 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n5 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t10 183.099
R731 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t10 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n4 183.099
R732 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n0 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t12 182.653
R733 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t13 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n3 182.297
R734 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n0 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t15 182.288
R735 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n7 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t6 182.285
R736 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n5 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t7 182.263
R737 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t6 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n6 182.263
R738 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t7 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n4 182.263
R739 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n20 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t2 155.667
R740 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n19 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t0 155.667
R741 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t11 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n2 146.282
R742 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n12 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t8 145.889
R743 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t8 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n11 145.857
R744 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n9 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t11 145.851
R745 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n14 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t5 135.911
R746 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n17 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n16 122.928
R747 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n20 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n19 109.715
R748 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t9 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n15 98.2234
R749 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n17 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t9 49.4098
R750 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n1 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t14 45.8204
R751 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n14 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n1 28.5785
R752 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n16 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t4 28.5685
R753 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t5 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n13 19.7637
R754 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n18 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n17 5.00095
R755 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n10 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n2 4.13208
R756 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n21 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t3 3.16453
R757 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n15 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n14 2.83669
R758 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n18 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n0 1.3453
R759 pmu_circuits_0.ring_100mV_0.mdls_inv_6.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n21 1.29092
R760 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n6 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n5 0.835457
R761 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n8 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n4 0.813812
R762 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n7 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n3 0.810242
R763 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n11 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n10 0.607643
R764 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n10 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n9 0.43198
R765 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n13 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN 0.339159
R766 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n12 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n2 0.333833
R767 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n9 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n8 0.21421
R768 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n11 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n3 0.21421
R769 pmu_circuits_0.ring_100mV_0.mdls_inv_6.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n18 0.184521
R770 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n12 0.120801
R771 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n8 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n7 0.106457
R772 gpio_analog[7].n7 gpio_analog[7].t7 206.963
R773 gpio_analog[7].n3 gpio_analog[7].t9 206.963
R774 gpio_analog[7].n3 gpio_analog[7].t5 206.321
R775 gpio_analog[7].n4 gpio_analog[7].t4 206.321
R776 gpio_analog[7].n5 gpio_analog[7].t0 206.321
R777 gpio_analog[7].n7 gpio_analog[7].t8 206.321
R778 gpio_analog[7].n9 gpio_analog[7].t6 206.321
R779 gpio_analog[7].n11 gpio_analog[7].t2 206.321
R780 gpio_analog[7].t5 gpio_analog[7].n2 206.317
R781 gpio_analog[7].t4 gpio_analog[7].n1 206.317
R782 gpio_analog[7].t0 gpio_analog[7].n0 206.317
R783 gpio_analog[7].t8 gpio_analog[7].n6 206.317
R784 gpio_analog[7].t6 gpio_analog[7].n8 206.317
R785 gpio_analog[7].t2 gpio_analog[7].n10 206.317
R786 pmu_circuits_0.ldo_iref gpio_analog[7] 187.281
R787 gpio_analog[7].n12 gpio_analog[7].t1 3.41293
R788 gpio_analog[7].n12 gpio_analog[7].t3 3.41293
R789 pmu_circuits_0.ldo_iref gpio_analog[7].n13 1.64033
R790 gpio_analog[7].n11 gpio_analog[7].n9 0.642396
R791 gpio_analog[7].n9 gpio_analog[7].n7 0.642396
R792 gpio_analog[7].n4 gpio_analog[7].n3 0.642396
R793 gpio_analog[7].n5 gpio_analog[7].n4 0.642396
R794 gpio_analog[7].n13 gpio_analog[7] 0.235123
R795 gpio_analog[7].n13 gpio_analog[7].n5 0.192876
R796 gpio_analog[7] gpio_analog[7].n12 0.184094
R797 gpio_analog[7].n13 gpio_analog[7].n11 0.183948
R798 a_350722_615130.n0 a_350722_615130.t0 7.40825
R799 a_350722_615130.n0 a_350722_615130.t3 4.70699
R800 a_350722_615130.n1 a_350722_615130.t4 4.53569
R801 a_350722_615130.t6 a_350722_615130.n5 4.53369
R802 a_350722_615130.n3 a_350722_615130.t7 4.38957
R803 a_350722_615130.n2 a_350722_615130.t5 4.3873
R804 a_350722_615130.n4 a_350722_615130.t1 4.26166
R805 a_350722_615130.n4 a_350722_615130.t2 4.06962
R806 a_350722_615130.n3 a_350722_615130.n2 2.26478
R807 a_350722_615130.n5 a_350722_615130.n4 2.0915
R808 a_350722_615130.n1 a_350722_615130.n0 0.66715
R809 a_350722_615130.n5 a_350722_615130.n3 0.1505
R810 a_350722_615130.n2 a_350722_615130.n1 0.144506
R811 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n2 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t0 265.382
R812 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n4 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n3 262.217
R813 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n10 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t5 183.099
R814 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n9 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t9 183.099
R815 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t9 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n8 183.099
R816 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n5 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t7 182.653
R817 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t5 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n0 182.297
R818 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n5 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t11 182.288
R819 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t8 182.285
R820 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n9 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t10 182.263
R821 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t8 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n10 182.263
R822 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t10 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n8 182.263
R823 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n2 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t4 155.667
R824 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n3 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t2 155.667
R825 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t12 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n7 146.282
R826 pmu_circuits_0.ring_100mV_0.mdls_inv_1.IN pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t6 145.889
R827 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t6 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n13 145.857
R828 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n11 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t12 145.851
R829 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n15 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t15 135.911
R830 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n18 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n17 122.928
R831 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n3 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n2 109.715
R832 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t13 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n16 98.2234
R833 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n18 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t13 49.4098
R834 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n6 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t14 45.8204
R835 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n15 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n6 28.5785
R836 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n17 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t1 28.5685
R837 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t15 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n14 19.7637
R838 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n16 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n15 5.198
R839 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n18 5.00095
R840 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n12 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n7 4.13208
R841 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n4 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t3 3.16453
R842 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n5 1.45868
R843 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n4 1.36143
R844 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n10 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n9 0.835457
R845 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n8 0.813812
R846 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n0 0.810242
R847 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n13 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n12 0.607643
R848 pmu_circuits_0.ring_100mV_0.mdls_inv_1.IN pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n7 0.454134
R849 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n12 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n11 0.43198
R850 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n14 pmu_circuits_0.ring_100mV_0.mdls_inv_1.IN 0.339159
R851 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n11 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n1 0.320167
R852 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n13 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n0 0.21421
R853 a_341818_613263.n1 a_341818_613263.t3 260.2
R854 a_341818_613263.n0 a_341818_613263.t6 252.136
R855 a_341818_613263.t5 a_341818_613263.n4 251.333
R856 a_341818_613263.n2 a_341818_613263.n0 164.748
R857 a_341818_613263.n4 a_341818_613263.t1 157.893
R858 a_341818_613263.n3 a_341818_613263.t4 155.667
R859 a_341818_613263.n1 a_341818_613263.t2 149.827
R860 a_341818_613263.n3 a_341818_613263.n2 72.9605
R861 a_341818_613263.n2 a_341818_613263.n1 9.14336
R862 a_341818_613263.n4 a_341818_613263.n3 8.74717
R863 a_341818_613263.n0 a_341818_613263.t0 3.16453
R864 a_345642_616040.t5 a_345642_616040.n4 260.2
R865 a_345642_616040.n2 a_345642_616040.t6 252.136
R866 a_345642_616040.n0 a_345642_616040.t4 251.333
R867 a_345642_616040.n3 a_345642_616040.n2 164.748
R868 a_345642_616040.n0 a_345642_616040.t1 157.893
R869 a_345642_616040.n1 a_345642_616040.t2 155.667
R870 a_345642_616040.n4 a_345642_616040.t3 149.827
R871 a_345642_616040.n3 a_345642_616040.n1 72.9605
R872 a_345642_616040.n4 a_345642_616040.n3 9.14336
R873 a_345642_616040.n1 a_345642_616040.n0 8.74717
R874 a_345642_616040.n2 a_345642_616040.t0 3.16453
R875 io_out[16].n1 io_out[16] 219.25
R876 io_out[16].n0 io_out[16].t1 147.147
R877 io_out[16].n0 io_out[16].t0 63.6678
R878 io_out[16] io_out[16].n0 44.5008
R879 pmu_circuits_0.ldo_vs io_out[16] 0.0700122
R880 io_out[16].n1 pmu_circuits_0.ldo_vs 0.0663537
R881 pmu_circuits_0.ldo_vs io_out[16].n1 0.061586
R882 io_out[15].n6 io_out[15].n5 4888.24
R883 io_out[15].n9 io_out[15].n6 4884.71
R884 io_out[15].n17 io_out[15].n4 1355.29
R885 io_out[15].n13 io_out[15].n11 1351.76
R886 io_out[15].n7 io_out[15].n3 521.413
R887 io_out[15].n8 io_out[15].n7 521.035
R888 io_out[15].n18 io_out[15].n3 376.848
R889 io_out[15].n8 io_out[15].n2 357.647
R890 io_out[15].n16 io_out[15].n15 271.43
R891 io_out[15].n14 io_out[15].n10 270.724
R892 io_out[15].n16 io_out[15].n5 261.185
R893 io_out[15].n10 io_out[15].n9 229.173
R894 io_out[15].n25 io_out[15] 199.394
R895 io_out[15].n20 io_out[15].n18 74.0415
R896 io_out[15].n20 io_out[15].n2 72.1843
R897 io_out[15].t0 io_out[15].n14 31.8085
R898 io_out[15].n1 io_out[15].t1 7.2144
R899 io_out[15].n24 io_out[15].t4 5.74557
R900 io_out[15].n19 io_out[15].t2 4.7068
R901 io_out[15].n20 io_out[15].n19 4.49173
R902 io_out[15].n15 io_out[15].t0 4.24157
R903 io_out[15].n21 io_out[15].n0 3.31278
R904 io_out[15].n21 io_out[15].n20 1.23559
R905 io_out[15].n24 io_out[15].t3 0.292821
R906 io_out[15].n24 io_out[15].n23 0.234051
R907 io_out[15] io_out[15].n24 0.216265
R908 pmu_circuits_0.ldo_out io_out[15] 0.124626
R909 io_out[15].n22 io_out[15].n1 0.0383289
R910 io_out[15].n23 io_out[15].n22 0.033381
R911 io_out[15].n25 pmu_circuits_0.ldo_out 0.0302203
R912 pmu_circuits_0.ldo_out io_out[15].n25 0.0257475
R913 io_out[15].n19 io_out[15].n1 0.0187887
R914 io_out[15].n11 io_out[15].n2 0.0153511
R915 io_out[15].n11 io_out[15].n10 0.014836
R916 io_out[15].n18 io_out[15].n17 0.0131168
R917 io_out[15].n17 io_out[15].n16 0.012684
R918 io_out[15].n12 io_out[15].n4 0.0069195
R919 io_out[15].n15 io_out[15].n4 0.00641981
R920 io_out[15].n13 io_out[15].n12 0.00449474
R921 io_out[15].n23 io_out[15].n0 0.00445473
R922 io_out[15].n5 io_out[15].n3 0.00432563
R923 io_out[15].n9 io_out[15].n8 0.00432563
R924 io_out[15].n14 io_out[15].n13 0.00399493
R925 io_out[15].n7 io_out[15].n6 0.00345991
R926 io_out[15].n15 io_out[15].n6 0.00345991
R927 io_out[15].n12 io_out[15].n0 0.00100012
R928 io_out[15].n22 io_out[15].n21 0.000504061
R929 a_352038_622652.n1 a_352038_622652.t0 177.476
R930 a_352038_622652.n2 a_352038_622652.t2 177.371
R931 a_352038_622652.n3 a_352038_622652.t6 31.4497
R932 a_352038_622652.n0 a_352038_622652.t4 17.6491
R933 a_352038_622652.n5 a_352038_622652.t5 10.2714
R934 a_352038_622652.n1 a_352038_622652.t1 4.93845
R935 a_352038_622652.t3 a_352038_622652.n0 2.90106
R936 a_352038_622652.n0 a_352038_622652.n3 0.941548
R937 a_352038_622652.n5 a_352038_622652.n4 0.923627
R938 a_352038_622652.n0 a_352038_622652.n7 0.836115
R939 a_352038_622652.n7 a_352038_622652.n6 0.773938
R940 a_352038_622652.n3 a_352038_622652.n2 0.288679
R941 a_352038_622652.n7 a_352038_622652.n5 0.224162
R942 a_352038_622652.n2 a_352038_622652.n1 0.0967847
R943 io_out[11].n4 io_out[11] 199.429
R944 io_out[11].n2 io_out[11].t1 21.3068
R945 io_out[11].n4 pmu_circuits_0.vref 18.0025
R946 io_out[11].n3 io_out[11].n1 11.9344
R947 io_out[11].n0 io_out[11].t2 11.7578
R948 io_out[11].n0 io_out[11].t3 11.7552
R949 io_out[11].n2 io_out[11].t0 10.1983
R950 pmu_circuits_0.iref io_out[11].n4 4.12586
R951 io_out[11].n3 io_out[11].n2 1.60834
R952 pmu_circuits_0.iref_2nA_0.IREF io_out[11] 1.46918
R953 io_out[11].n1 io_out[11].t4 1.05273
R954 pmu_circuits_0.vref io_out[11].n3 0.979689
R955 io_out[11] io_out[11].n0 0.151738
R956 pmu_circuits_0.iref pmu_circuits_0.iref_2nA_0.IREF 0.0540699
R957 io_out[11].n1 pmu_circuits_0.vref01_0.VREF 0.0165714
R958 a_341818_619927.n4 a_341818_619927.t3 260.2
R959 a_341818_619927.n2 a_341818_619927.t6 252.136
R960 a_341818_619927.n0 a_341818_619927.t2 251.333
R961 a_341818_619927.n3 a_341818_619927.n2 164.748
R962 a_341818_619927.n0 a_341818_619927.t1 157.893
R963 a_341818_619927.n1 a_341818_619927.t4 155.667
R964 a_341818_619927.t5 a_341818_619927.n4 149.827
R965 a_341818_619927.n3 a_341818_619927.n1 72.9605
R966 a_341818_619927.n4 a_341818_619927.n3 9.14336
R967 a_341818_619927.n1 a_341818_619927.n0 8.74717
R968 a_341818_619927.n2 a_341818_619927.t0 3.16453
R969 a_345642_617706.n0 a_345642_617706.t1 260.2
R970 a_345642_617706.n1 a_345642_617706.t6 252.136
R971 a_345642_617706.t3 a_345642_617706.n4 251.333
R972 a_345642_617706.n2 a_345642_617706.n1 164.748
R973 a_345642_617706.n4 a_345642_617706.t4 157.893
R974 a_345642_617706.n3 a_345642_617706.t2 155.667
R975 a_345642_617706.n0 a_345642_617706.t0 149.827
R976 a_345642_617706.n3 a_345642_617706.n2 72.9605
R977 a_345642_617706.n2 a_345642_617706.n0 9.14336
R978 a_345642_617706.n4 a_345642_617706.n3 8.74717
R979 a_345642_617706.n1 a_345642_617706.t5 3.16453
R980 a_335719_622037.n0 a_335719_622037.n6 113.371
R981 a_335719_622037.n5 a_335719_622037.n4 113.371
R982 a_335719_622037.n7 a_335719_622037.t9 74.6407
R983 a_335719_622037.n2 a_335719_622037.t8 74.6407
R984 a_335719_622037.t0 a_335719_622037.n3 73.5102
R985 a_335719_622037.t2 a_335719_622037.n8 73.5102
R986 a_335719_622037.n4 a_335719_622037.t7 73.5085
R987 a_335719_622037.n0 a_335719_622037.t2 73.5085
R988 a_335719_622037.n6 a_335719_622037.t6 73.5085
R989 a_335719_622037.n5 a_335719_622037.t0 73.5085
R990 a_335719_622037.n1 a_335719_622037.t5 14.0533
R991 a_335719_622037.n1 a_335719_622037.t4 11.7371
R992 a_335719_622037.t3 a_335719_622037.n0 7.79415
R993 a_335719_622037.n0 a_335719_622037.t1 7.49661
R994 a_335719_622037.n0 a_335719_622037.n1 5.59997
R995 a_335719_622037.n8 a_335719_622037.n7 1.13093
R996 a_335719_622037.n3 a_335719_622037.n2 1.13093
R997 a_335719_622037.n0 a_335719_622037.n5 0.985754
R998 a_341818_618261.n1 a_341818_618261.t2 260.2
R999 a_341818_618261.n0 a_341818_618261.t0 252.136
R1000 a_341818_618261.n3 a_341818_618261.t1 251.333
R1001 a_341818_618261.n2 a_341818_618261.n0 164.748
R1002 a_341818_618261.n3 a_341818_618261.t6 157.893
R1003 a_341818_618261.t4 a_341818_618261.n4 155.667
R1004 a_341818_618261.n1 a_341818_618261.t3 149.827
R1005 a_341818_618261.n4 a_341818_618261.n2 72.9605
R1006 a_341818_618261.n2 a_341818_618261.n1 9.14336
R1007 a_341818_618261.n4 a_341818_618261.n3 8.74717
R1008 a_341818_618261.n0 a_341818_618261.t5 3.16453
R1009 a_336843_616061.n0 a_336843_616061.t0 57.4135
R1010 a_336843_616061.n0 a_336843_616061.t2 9.98238
R1011 a_336843_616061.t1 a_336843_616061.n0 9.18355
R1012 a_345642_621038.n4 a_345642_621038.t3 260.2
R1013 a_345642_621038.n2 a_345642_621038.t6 252.136
R1014 a_345642_621038.n0 a_345642_621038.t2 251.333
R1015 a_345642_621038.n3 a_345642_621038.n2 164.748
R1016 a_345642_621038.n0 a_345642_621038.t1 157.893
R1017 a_345642_621038.n1 a_345642_621038.t4 155.667
R1018 a_345642_621038.t5 a_345642_621038.n4 149.827
R1019 a_345642_621038.n3 a_345642_621038.n1 72.9605
R1020 a_345642_621038.n4 a_345642_621038.n3 9.14336
R1021 a_345642_621038.n1 a_345642_621038.n0 8.74717
R1022 a_345642_621038.n2 a_345642_621038.t0 3.16453
R1023 a_345642_619372.n0 a_345642_619372.t1 260.2
R1024 a_345642_619372.n1 a_345642_619372.t0 252.136
R1025 a_345642_619372.t4 a_345642_619372.n4 251.333
R1026 a_345642_619372.n2 a_345642_619372.n1 164.748
R1027 a_345642_619372.n4 a_345642_619372.t5 157.893
R1028 a_345642_619372.n3 a_345642_619372.t3 155.667
R1029 a_345642_619372.n0 a_345642_619372.t2 149.827
R1030 a_345642_619372.n3 a_345642_619372.n2 72.9605
R1031 a_345642_619372.n2 a_345642_619372.n0 9.14336
R1032 a_345642_619372.n4 a_345642_619372.n3 8.74717
R1033 a_345642_619372.n1 a_345642_619372.t6 3.16453
R1034 a_345642_614374.n0 a_345642_614374.t4 260.2
R1035 a_345642_614374.n1 a_345642_614374.t0 252.136
R1036 a_345642_614374.n3 a_345642_614374.t6 251.333
R1037 a_345642_614374.n2 a_345642_614374.n1 164.748
R1038 a_345642_614374.n3 a_345642_614374.t1 157.893
R1039 a_345642_614374.t5 a_345642_614374.n4 155.667
R1040 a_345642_614374.n0 a_345642_614374.t3 149.827
R1041 a_345642_614374.n4 a_345642_614374.n2 72.9605
R1042 a_345642_614374.n2 a_345642_614374.n0 9.14336
R1043 a_345642_614374.n4 a_345642_614374.n3 8.74717
R1044 a_345642_614374.n1 a_345642_614374.t2 3.16453
R1045 pmu_circuits_0.ldo_vb io_out[12] 195.081
R1046 io_out[12].n0 io_out[12].t1 49.9518
R1047 io_out[12].n0 io_out[12].t0 48.1905
R1048 io_out[12] io_out[12].n0 2.75644
R1049 pmu_circuits_0.ldo_vb io_out[12] 0.0847338
C0 io_in[4] io_in_3v3[4] 0.0824f
C1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT 1.52f
C2 la_oenb[106] la_data_out[106] 0.0566f
C3 la_oenb[82] la_data_in[83] 0.0566f
C4 la_data_out[5] la_oenb[5] 0.0566f
C5 io_out[3] io_in[3] 0.0824f
C6 wbs_ack_o wbs_cyc_i 0.0566f
C7 io_out[12] io_out[15] 2.34f
C8 la_data_out[97] la_data_in[97] 0.0566f
C9 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN 0.0308f
C10 wbs_dat_o[10] wbs_adr_i[11] 0.0566f
C11 la_oenb[124] la_data_in[125] 0.0566f
C12 la_data_in[66] la_data_out[66] 0.0566f
C13 gpio_noesd[2] io_in_3v3[9] 0.0824f
C14 la_data_in[95] la_data_out[95] 0.0566f
C15 la_data_in[34] la_data_out[34] 0.0566f
C16 la_data_out[83] la_data_in[83] 0.0566f
C17 la_oenb[5] la_data_in[6] 0.0566f
C18 la_data_out[115] la_oenb[115] 0.0566f
C19 gpio_analog[12] gpio_noesd[12] 0.0824f
C20 gpio_noesd[6] gpio_analog[6] 0.0824f
C21 io_oeb[2] io_in_3v3[3] 0.0824f
C22 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_343294_617413# 6.45e-19
C23 io_in[9] io_in_3v3[9] 0.0824f
C24 la_data_in[90] la_data_out[90] 0.0566f
C25 io_clamp_high[0] io_analog[4] 1.2f
C26 la_data_out[9] la_oenb[9] 0.0566f
C27 la_oenb[125] la_data_in[126] 0.0566f
C28 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1 1.14f
C29 io_out[12] gpio_analog[3] 13.4f
C30 la_oenb[112] la_data_in[113] 0.0566f
C31 wbs_adr_i[31] wbs_dat_i[31] 0.0566f
C32 wbs_dat_i[28] wbs_dat_o[28] 0.0566f
C33 wbs_dat_o[29] wbs_adr_i[30] 0.0566f
C34 la_data_in[6] la_data_out[6] 0.0566f
C35 la_data_in[65] la_data_out[65] 0.0566f
C36 la_data_in[104] la_data_out[104] 0.0566f
C37 wbs_adr_i[24] wbs_dat_i[24] 0.0566f
C38 wbs_dat_i[1] wbs_dat_o[1] 0.0566f
C39 a_337674_621712# a_337674_622496# 1.17f
C40 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT io_out[12] 6.11e-19
C41 la_data_out[99] la_oenb[99] 0.0566f
C42 la_data_out[81] la_data_in[81] 0.0566f
C43 la_oenb[22] la_data_in[23] 0.0566f
C44 a_337674_621712# pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.00384f
C45 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT vccd1 0.144f
C46 wbs_dat_o[20] wbs_dat_i[20] 0.0566f
C47 wbs_dat_o[12] wbs_dat_i[12] 0.0566f
C48 la_data_out[61] la_data_in[61] 0.0566f
C49 la_data_out[70] la_oenb[70] 0.0566f
C50 io_in[14] io_out[14] 0.0824f
C51 a_345642_618736# pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT 1.09f
C52 io_in_3v3[11] io_in[11] 0.0824f
C53 a_345642_615404# pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT 0.00146f
C54 wbs_adr_i[26] wbs_dat_o[25] 0.0566f
C55 wbs_cyc_i wbs_stb_i 0.0566f
C56 io_out[11] pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 1.16f
C57 io_out[16] io_out[12] 1.02f
C58 wbs_adr_i[18] wbs_dat_o[17] 0.0566f
C59 io_clamp_low[0] io_clamp_high[0] 0.711f
C60 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT 1.75f
C61 la_data_in[42] la_data_out[42] 0.0566f
C62 wbs_dat_i[19] wbs_dat_o[19] 0.0566f
C63 la_data_out[115] la_data_in[115] 0.0566f
C64 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 9.45e-20
C65 la_oenb[12] la_data_out[12] 0.0566f
C66 la_data_out[89] la_oenb[89] 0.0566f
C67 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT 0.112f
C68 io_in[7] io_in_3v3[7] 0.0824f
C69 la_oenb[110] la_data_out[110] 0.0566f
C70 la_oenb[34] la_data_in[35] 0.0566f
C71 a_337674_622496# pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg 0.156f
C72 la_data_out[109] la_oenb[109] 0.0566f
C73 la_data_in[71] la_data_out[71] 0.0566f
C74 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN vccd1 0.172f
C75 m3_583220_500050# io_out[12] 0.00631f
C76 la_data_out[93] la_data_in[93] 0.0566f
C77 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.354f
C78 wbs_dat_o[8] wbs_adr_i[9] 0.0566f
C79 io_out[16] io_in[16] 0.0824f
C80 la_data_out[119] la_data_in[119] 0.0566f
C81 la_data_out[79] la_oenb[79] 0.0566f
C82 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT 4.97f
C83 la_data_out[60] la_oenb[60] 0.0566f
C84 io_oeb[4] io_out[4] 0.0824f
C85 la_data_out[125] la_data_in[125] 0.0566f
C86 io_out[4] io_in[4] 0.0824f
C87 la_oenb[75] la_data_in[76] 0.0566f
C88 m3_326794_701100# io_analog[4] 0.00974f
C89 a_345642_613738# pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT 1.21f
C90 wbs_adr_i[11] wbs_dat_i[11] 0.0566f
C91 la_data_in[36] la_data_out[36] 0.0566f
C92 a_337674_621712# vccd1 0.784f
C93 w_336471_617254# a_336716_619863# 6.92e-21
C94 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT io_out[11] 0.963f
C95 wbs_adr_i[17] wbs_dat_i[17] 0.0566f
C96 wbs_stb_i wbs_we_i 0.0566f
C97 la_oenb[72] la_data_out[72] 0.0566f
C98 wbs_adr_i[15] wbs_dat_i[15] 0.0566f
C99 la_oenb[47] la_data_in[48] 0.0566f
C100 la_data_in[54] la_data_out[54] 0.0566f
C101 la_data_in[103] la_data_out[103] 0.0566f
C102 io_in_3v3[26] io_in[26] 0.0824f
C103 la_data_out[105] la_oenb[105] 0.0566f
C104 vssd1 io_out[11] 2.84f
C105 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT 2.35f
C106 vccd1 io_out[11] 5.81f
C107 io_in_3v3[13] io_in[13] 0.0824f
C108 la_data_out[85] la_oenb[85] 0.0566f
C109 la_oenb[60] la_data_in[61] 0.0566f
C110 la_oenb[114] la_data_in[115] 0.0566f
C111 la_data_out[6] la_oenb[6] 0.0566f
C112 io_in[6] io_in_3v3[6] 0.0824f
C113 io_clamp_low[1] io_analog[5] 0.972f
C114 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_345642_615404# 0.876f
C115 a_343294_620745# pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN 1.37e-19
C116 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_343294_619079# 1.08f
C117 la_data_out[117] la_oenb[117] 0.0566f
C118 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN vccd1 0.0999f
C119 io_out[18] io_in[18] 0.0824f
C120 wbs_dat_i[13] wbs_dat_o[13] 0.0566f
C121 la_oenb[46] la_data_in[47] 0.0566f
C122 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT 0.121f
C123 a_343294_617413# vdda1 1.59f
C124 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT 0.192f
C125 io_out[1] io_in[1] 0.0824f
C126 io_oeb[11] io_out[11] 0.0968f
C127 la_oenb[42] la_data_in[43] 0.0566f
C128 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 7.84e-20
C129 la_data_out[88] la_oenb[88] 0.0566f
C130 m3_326794_701100# io_clamp_low[0] 0.00389f
C131 a_339370_617808# pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.361f
C132 la_oenb[83] la_data_in[84] 0.0566f
C133 vccd1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg 0.51f
C134 wbs_adr_i[8] wbs_dat_i[8] 0.0566f
C135 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1 a_336716_619863# 0.595f
C136 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN 1.46f
C137 vdda1 a_343294_619079# 1.59f
C138 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT 0.179f
C139 vccd1 vdda1 1.73f
C140 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_345642_617070# 1.22f
C141 la_data_in[21] la_data_out[21] 0.0566f
C142 la_data_in[124] la_data_out[124] 0.0566f
C143 io_in[8] io_out[8] 0.0824f
C144 la_data_in[108] la_data_out[108] 0.0566f
C145 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_345642_615404# 1.09f
C146 gpio_noesd[1] gpio_analog[1] 0.0824f
C147 io_oeb[13] io_out[13] 0.0824f
C148 wbs_adr_i[21] wbs_dat_i[21] 0.0566f
C149 io_in[15] io_in_3v3[15] 0.0824f
C150 gpio_noesd[9] io_in_3v3[16] 0.0824f
C151 la_data_in[18] la_oenb[17] 0.0566f
C152 la_data_out[1] la_oenb[1] 0.0566f
C153 la_data_out[1] la_data_in[1] 0.0566f
C154 wbs_adr_i[6] wbs_dat_i[6] 0.0566f
C155 wbs_dat_i[5] wbs_dat_o[5] 0.0566f
C156 la_data_in[28] la_data_out[28] 0.0566f
C157 wbs_dat_o[5] wbs_adr_i[6] 0.0566f
C158 la_data_out[111] la_data_in[111] 0.0566f
C159 wbs_adr_i[24] wbs_dat_o[23] 0.0566f
C160 la_data_in[112] la_data_out[112] 0.0566f
C161 la_oenb[107] la_data_in[108] 0.0566f
C162 la_data_out[11] la_oenb[11] 0.0566f
C163 io_in_3v3[8] gpio_noesd[1] 0.0824f
C164 la_data_in[46] la_data_out[46] 0.0566f
C165 la_data_out[125] la_oenb[125] 0.0566f
C166 la_data_out[49] la_oenb[49] 0.0566f
C167 la_oenb[98] la_data_out[98] 0.0566f
C168 gpio_noesd[12] io_in_3v3[19] 0.0824f
C169 m3_222594_700786# m3_225094_700796# 0.00779f
C170 la_data_in[117] la_data_out[117] 0.0566f
C171 wbs_dat_i[11] wbs_dat_o[11] 0.0566f
C172 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT 4.71f
C173 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT a_339370_617808# 3.09e-19
C174 la_oenb[55] la_data_in[56] 0.0566f
C175 la_data_out[107] la_oenb[107] 0.0566f
C176 wbs_dat_o[6] wbs_dat_i[6] 0.0566f
C177 vccd1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT 0.00217f
C178 la_data_in[116] la_oenb[115] 0.0566f
C179 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_345642_617070# 6.99e-19
C180 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT a_343294_614081# 0.607f
C181 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT 0.0308f
C182 vccd1 a_339370_617808# 0.709f
C183 io_in_3v3[2] io_in[2] 0.0824f
C184 io_in_3v3[7] gpio_noesd[0] 0.0824f
C185 la_data_in[91] la_data_out[91] 0.0566f
C186 io_in[7] io_out[7] 0.0824f
C187 la_oenb[90] la_data_in[91] 0.0566f
C188 io_in_3v3[20] gpio_noesd[13] 0.0824f
C189 io_in[10] io_in_3v3[10] 0.0824f
C190 la_data_in[88] la_data_out[88] 0.0566f
C191 la_data_in[82] la_data_out[82] 0.0566f
C192 la_oenb[85] la_data_in[86] 0.0566f
C193 la_data_in[47] la_data_out[47] 0.0566f
C194 io_oeb[6] io_out[6] 0.0824f
C195 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 a_336716_619863# 0.32f
C196 la_data_in[12] la_oenb[11] 0.0566f
C197 a_345642_618736# pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN 0.00146f
C198 la_oenb[126] la_data_in[127] 0.0566f
C199 io_out[6] io_in[6] 0.0824f
C200 la_oenb[1] la_data_in[2] 0.0566f
C201 user_irq[1] user_irq[0] 0.0566f
C202 wbs_dat_o[6] wbs_adr_i[7] 0.0566f
C203 la_oenb[102] la_data_out[102] 0.0566f
C204 la_oenb[63] la_data_in[64] 0.0566f
C205 la_oenb[118] la_data_in[119] 0.0566f
C206 la_data_out[89] la_data_in[89] 0.0566f
C207 la_data_out[107] la_data_in[107] 0.0566f
C208 la_oenb[28] la_data_in[29] 0.0566f
C209 gpio_analog[7] io_out[15] 9.67f
C210 la_data_in[23] la_data_out[23] 0.0566f
C211 la_data_in[85] la_data_out[85] 0.0566f
C212 wbs_adr_i[8] wbs_dat_o[7] 0.0566f
C213 io_in_3v3[1] io_oeb[0] 0.0824f
C214 wbs_adr_i[18] wbs_dat_i[18] 0.0566f
C215 la_oenb[40] la_data_in[41] 0.0566f
C216 la_data_in[72] la_data_out[72] 0.0566f
C217 io_out[23] io_oeb[23] 0.0824f
C218 la_data_in[80] la_data_out[80] 0.0566f
C219 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT 2.12f
C220 la_oenb[119] la_data_in[120] 0.0566f
C221 io_oeb[7] io_out[7] 0.0824f
C222 la_oenb[58] la_data_in[59] 0.0566f
C223 la_data_in[13] la_data_out[13] 0.0566f
C224 wbs_adr_i[22] wbs_dat_i[22] 0.0566f
C225 gpio_noesd[7] io_in_3v3[14] 0.0824f
C226 a_345642_615404# vdda1 1.59f
C227 io_in[5] io_in_3v3[5] 0.0824f
C228 wbs_dat_i[29] wbs_dat_o[29] 0.0566f
C229 la_oenb[54] la_data_in[55] 0.0566f
C230 la_oenb[29] la_data_in[30] 0.0566f
C231 la_oenb[23] la_data_in[24] 0.0566f
C232 la_data_in[110] la_data_out[110] 0.0566f
C233 m3_170894_700738# m3_173394_700736# 0.00935f
C234 la_data_in[12] la_data_out[12] 0.0566f
C235 la_data_out[42] la_oenb[42] 0.0566f
C236 la_data_out[45] la_data_in[45] 0.0566f
C237 wbs_dat_i[15] wbs_dat_o[15] 0.0566f
C238 la_data_in[17] la_data_out[17] 0.0566f
C239 la_oenb[106] la_data_in[107] 0.0566f
C240 la_data_in[28] la_oenb[27] 0.0566f
C241 la_data_out[82] la_oenb[82] 0.0566f
C242 la_oenb[116] la_data_in[117] 0.0566f
C243 la_data_in[57] la_data_out[57] 0.0566f
C244 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_345642_613738# 1.29e-19
C245 io_out[11] a_339370_618592# 0.157f
C246 la_data_in[2] la_data_out[2] 0.0566f
C247 la_data_out[35] la_data_in[35] 0.0566f
C248 wbs_dat_i[7] wbs_adr_i[7] 0.0566f
C249 la_oenb[90] la_data_out[90] 0.0566f
C250 la_oenb[50] la_data_in[51] 0.0566f
C251 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_345642_620402# 0.603f
C252 vssd1 io_out[15] 1.12f
C253 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT a_336716_619863# 0.264f
C254 la_data_in[9] la_data_out[9] 0.0566f
C255 vccd1 io_out[15] 2.23f
C256 wbs_dat_o[14] wbs_dat_i[14] 0.0566f
C257 wbs_we_i wbs_adr_i[0] 0.0566f
C258 la_data_in[58] la_data_out[58] 0.0566f
C259 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_343294_617413# 0.00194f
C260 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT 2.12f
C261 wbs_dat_i[24] wbs_dat_o[24] 0.0566f
C262 vccd1 a_336716_619863# 0.00177f
C263 gpio_analog[7] io_out[16] 0.00227f
C264 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT 4.57f
C265 a_345642_617070# vdda1 1.59f
C266 la_data_in[98] la_data_out[98] 0.0566f
C267 la_oenb[53] la_data_in[54] 0.0566f
C268 la_data_out[61] la_oenb[61] 0.0566f
C269 wbs_adr_i[10] wbs_dat_o[9] 0.0566f
C270 io_oeb[24] io_in_3v3[25] 0.0824f
C271 la_data_out[13] la_oenb[13] 0.0566f
C272 la_oenb[44] la_data_in[45] 0.0566f
C273 la_data_in[104] la_oenb[103] 0.0566f
C274 wbs_dat_o[0] wbs_dat_i[0] 0.0566f
C275 la_data_in[114] la_oenb[113] 0.0566f
C276 io_in_3v3[18] io_in[18] 0.0824f
C277 la_data_in[0] la_data_out[0] 0.0566f
C278 vssd1 gpio_analog[3] 2.23f
C279 vccd1 gpio_analog[3] 4.28f
C280 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT a_343294_615747# 2.93e-21
C281 a_343294_614081# pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT 1.07f
C282 la_data_out[94] la_oenb[94] 0.0566f
C283 la_oenb[73] la_data_in[74] 0.0566f
C284 m3_583180_455628# io_out[11] 0.00746f
C285 io_in_3v3[23] gpio_noesd[16] 0.0824f
C286 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_343294_619079# 0.00136f
C287 a_345642_620402# vdda1 1.59f
C288 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT vccd1 0.144f
C289 la_data_out[3] la_data_in[3] 0.0566f
C290 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_345642_613738# 0.669f
C291 io_out[1] io_oeb[1] 0.0824f
C292 la_data_out[104] la_oenb[104] 0.0566f
C293 la_data_in[53] la_data_out[53] 0.0566f
C294 wbs_dat_i[7] wbs_dat_o[7] 0.0566f
C295 io_in_3v3[18] gpio_noesd[11] 0.0824f
C296 wbs_dat_o[11] wbs_adr_i[12] 0.0566f
C297 la_data_out[15] la_oenb[15] 0.0566f
C298 la_oenb[46] la_data_out[46] 0.0566f
C299 la_data_out[37] la_oenb[37] 0.0566f
C300 la_data_in[86] la_data_out[86] 0.0566f
C301 io_out[19] io_oeb[19] 0.0824f
C302 la_data_out[39] la_oenb[39] 0.0566f
C303 la_oenb[100] la_data_out[100] 0.0566f
C304 la_data_in[26] la_data_out[26] 0.0566f
C305 io_out[17] io_oeb[17] 0.0824f
C306 vssd1 io_out[16] 3.63f
C307 io_out[16] vccd1 0.874f
C308 la_data_in[43] la_data_out[43] 0.0566f
C309 la_oenb[41] la_data_in[42] 0.0566f
C310 io_in_3v3[11] gpio_noesd[4] 0.0824f
C311 io_in[11] io_out[11] 0.0824f
C312 wbs_dat_o[16] wbs_adr_i[17] 0.0566f
C313 io_in_3v3[22] io_in[22] 0.0824f
C314 la_data_in[94] la_oenb[93] 0.0566f
C315 la_data_out[54] la_oenb[54] 0.0566f
C316 gpio_analog[11] gpio_noesd[11] 0.0824f
C317 wbs_dat_i[23] wbs_dat_o[23] 0.0566f
C318 la_data_out[27] la_oenb[27] 0.0566f
C319 la_data_out[83] la_oenb[83] 0.0566f
C320 wbs_dat_i[5] wbs_adr_i[5] 0.0566f
C321 gpio_analog[15] gpio_noesd[15] 0.0824f
C322 io_out[17] io_in[17] 0.0824f
C323 la_data_out[96] la_oenb[96] 0.0566f
C324 la_data_out[101] la_oenb[101] 0.0566f
C325 la_oenb[68] la_data_in[69] 0.0566f
C326 la_oenb[9] la_data_in[10] 0.0566f
C327 a_345642_615404# a_343294_615747# 0.0129f
C328 io_clamp_low[0] io_analog[4] 1.2f
C329 la_data_out[29] la_data_in[29] 0.0566f
C330 la_oenb[76] la_data_in[77] 0.0566f
C331 wbs_dat_i[22] wbs_dat_o[22] 0.0566f
C332 la_data_in[105] la_data_out[105] 0.0566f
C333 la_data_out[79] la_data_in[79] 0.0566f
C334 io_out[5] io_in[5] 0.0824f
C335 la_oenb[15] la_data_in[16] 0.0566f
C336 a_339370_618592# a_339370_617808# 1.17f
C337 io_oeb[5] io_out[5] 0.0824f
C338 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT vdda1 4.65f
C339 a_343294_620745# pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT 6.45e-19
C340 la_data_out[28] la_oenb[28] 0.0566f
C341 la_oenb[14] la_data_in[15] 0.0566f
C342 la_data_in[127] la_data_out[127] 0.0566f
C343 la_data_in[87] la_data_out[87] 0.0566f
C344 io_in_3v3[19] io_in[19] 0.0824f
C345 wbs_dat_i[27] wbs_dat_o[27] 0.0566f
C346 wbs_dat_o[10] wbs_dat_i[10] 0.0566f
C347 io_out[20] io_oeb[20] 0.0824f
C348 la_oenb[16] la_data_in[17] 0.0566f
C349 la_oenb[69] la_data_in[70] 0.0566f
C350 la_data_in[19] la_data_out[19] 0.0566f
C351 la_data_out[33] la_oenb[33] 0.0566f
C352 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT a_343294_615747# 0.827f
C353 io_in[12] io_in_3v3[12] 0.0824f
C354 a_345642_613738# vdda1 1.59f
C355 la_oenb[56] la_data_in[57] 0.0566f
C356 io_out[18] io_oeb[18] 0.0824f
C357 la_data_out[118] la_oenb[118] 0.0566f
C358 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_345642_615404# 1.06e-19
C359 gpio_noesd[4] gpio_analog[4] 0.0824f
C360 la_data_in[116] la_data_out[116] 0.0566f
C361 la_oenb[18] la_data_in[19] 0.0566f
C362 la_data_in[16] la_data_out[16] 0.0566f
C363 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 1.03e-19
C364 io_oeb[26] io_out[26] 0.0824f
C365 a_345642_613738# a_343294_614081# 0.0129f
C366 la_oenb[94] la_data_in[95] 0.0566f
C367 la_oenb[127] user_clock2 0.0566f
C368 wbs_adr_i[4] wbs_dat_i[4] 0.0566f
C369 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN vdda1 4.59f
C370 io_in_3v3[10] gpio_noesd[3] 0.0824f
C371 a_337674_621712# pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg 0.011f
C372 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT 0.179f
C373 la_data_out[51] la_oenb[51] 0.0566f
C374 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_343294_614081# 0.00194f
C375 la_data_in[40] la_oenb[39] 0.0566f
C376 la_data_out[24] la_oenb[24] 0.0566f
C377 wb_clk_i wb_rst_i 0.0566f
C378 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 1.23e-19
C379 la_oenb[38] la_data_out[38] 0.0566f
C380 wbs_dat_o[31] la_data_in[0] 0.0566f
C381 wbs_adr_i[16] wbs_dat_o[15] 0.0566f
C382 gpio_noesd[2] gpio_analog[2] 0.0824f
C383 wbs_dat_o[18] wbs_dat_i[18] 0.0566f
C384 la_data_in[37] la_data_out[37] 0.0566f
C385 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg io_out[11] 0.0774f
C386 la_oenb[97] la_data_in[98] 0.0566f
C387 la_oenb[123] la_data_in[124] 0.0566f
C388 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_345642_617070# 0.664f
C389 wbs_adr_i[20] wbs_dat_i[20] 0.0566f
C390 wbs_adr_i[26] wbs_dat_i[26] 0.0566f
C391 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN a_343294_617413# 0.664f
C392 wbs_adr_i[12] wbs_dat_i[12] 0.0566f
C393 vdda1 io_out[11] 4.81f
C394 m3_660_462398# io_out[15] 0.00772f
C395 la_data_out[75] la_data_in[75] 0.0566f
C396 la_data_out[31] la_oenb[31] 0.0566f
C397 la_oenb[81] la_data_in[82] 0.0566f
C398 wbs_adr_i[28] wbs_dat_i[28] 0.0566f
C399 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT a_345642_620402# 0.00215f
C400 wbs_dat_o[30] wbs_adr_i[31] 0.0566f
C401 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN vdda1 6.24f
C402 la_data_out[17] la_oenb[17] 0.0566f
C403 la_data_out[57] la_oenb[57] 0.0566f
C404 la_data_out[77] la_data_in[77] 0.0566f
C405 a_343294_617413# pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN 1.07f
C406 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN a_343294_619079# 3.18e-19
C407 wbs_dat_i[16] wbs_dat_o[16] 0.0566f
C408 la_data_in[44] la_data_out[44] 0.0566f
C409 a_345642_618736# pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT 0.876f
C410 la_oenb[26] la_data_in[27] 0.0566f
C411 wbs_dat_o[22] wbs_adr_i[23] 0.0566f
C412 io_clamp_low[2] io_clamp_high[2] 0.781f
C413 la_data_out[3] la_oenb[3] 0.0566f
C414 la_oenb[49] la_data_in[50] 0.0566f
C415 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN vccd1 0.0297f
C416 la_data_out[53] la_oenb[53] 0.0566f
C417 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT a_343294_615747# 0.00155f
C418 io_in[15] io_out[15] 0.0824f
C419 gpio_analog[13] gpio_noesd[13] 0.0824f
C420 la_oenb[2] la_data_in[3] 0.0566f
C421 wbs_adr_i[22] wbs_dat_o[21] 0.0566f
C422 io_out[9] io_in[9] 0.0824f
C423 la_oenb[30] la_data_in[31] 0.0566f
C424 gpio_analog[7] io_out[12] 0.454f
C425 la_data_in[38] la_oenb[37] 0.0566f
C426 la_data_out[111] la_oenb[111] 0.0566f
C427 la_oenb[52] la_data_in[53] 0.0566f
C428 la_data_in[78] la_data_out[78] 0.0566f
C429 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN a_343294_619079# 0.829f
C430 io_clamp_low[1] io_clamp_high[1] 0.77f
C431 user_irq[1] user_irq[2] 0.0566f
C432 vccd1 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN 0.0236f
C433 la_data_in[76] la_data_out[76] 0.0566f
C434 wbs_dat_o[1] wbs_sel_i[1] 0.0566f
C435 io_out[11] a_339370_617808# 0.00626f
C436 la_data_in[52] la_data_out[52] 0.0566f
C437 la_oenb[64] la_data_in[65] 0.0566f
C438 la_oenb[66] la_data_in[67] 0.0566f
C439 la_oenb[0] la_data_in[1] 0.0566f
C440 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT 1.46f
C441 io_in[26] io_out[26] 0.0824f
C442 vdda1 a_343294_614081# 1.59f
C443 wbs_dat_o[4] wbs_adr_i[5] 0.0566f
C444 gpio_analog[10] gpio_noesd[10] 0.0824f
C445 la_oenb[86] la_data_in[87] 0.0566f
C446 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN a_343294_615747# 0.00136f
C447 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT 2.1f
C448 la_oenb[126] la_data_out[126] 0.0566f
C449 la_data_in[40] la_data_out[40] 0.0566f
C450 la_oenb[12] la_data_in[13] 0.0566f
C451 vssd1 io_out[12] 2.84f
C452 io_out[12] vccd1 4.35f
C453 la_data_out[67] la_data_in[67] 0.0566f
C454 la_data_in[90] la_oenb[89] 0.0566f
C455 la_data_out[127] la_oenb[127] 0.0566f
C456 la_data_out[91] la_oenb[91] 0.0566f
C457 wbs_adr_i[1] wbs_dat_i[1] 0.0566f
C458 a_345642_618736# a_343294_619079# 0.0129f
C459 la_data_out[121] la_oenb[121] 0.0566f
C460 la_data_out[2] la_oenb[2] 0.0566f
C461 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT 4.8f
C462 gpio_analog[17] gpio_noesd[17] 0.0824f
C463 m3_326794_701100# m3_324294_701080# 0.00584f
C464 la_data_in[120] la_data_out[120] 0.0566f
C465 la_data_out[40] la_oenb[40] 0.0566f
C466 la_data_in[101] la_data_out[101] 0.0566f
C467 la_oenb[44] la_data_out[44] 0.0566f
C468 la_oenb[25] la_data_in[26] 0.0566f
C469 la_oenb[74] la_data_in[75] 0.0566f
C470 io_in[24] io_out[24] 0.0824f
C471 wbs_adr_i[3] wbs_dat_i[3] 0.0566f
C472 wbs_dat_o[24] wbs_adr_i[25] 0.0566f
C473 la_oenb[61] la_data_in[62] 0.0566f
C474 la_data_out[45] la_oenb[45] 0.0566f
C475 la_data_in[8] la_data_out[8] 0.0566f
C476 io_out[22] io_oeb[22] 0.0824f
C477 w_336471_617254# pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.118f
C478 io_in[21] io_out[21] 0.0824f
C479 la_data_out[26] la_oenb[26] 0.0566f
C480 la_oenb[16] la_data_out[16] 0.0566f
C481 wbs_dat_i[31] wbs_dat_o[31] 0.0566f
C482 io_out[10] io_in[10] 0.0824f
C483 la_data_in[48] la_data_out[48] 0.0566f
C484 la_data_out[0] la_oenb[0] 0.0566f
C485 la_data_out[87] la_oenb[87] 0.0566f
C486 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT 0.134f
C487 la_data_in[68] la_data_out[68] 0.0566f
C488 la_data_out[103] la_oenb[103] 0.0566f
C489 la_data_out[121] la_data_in[121] 0.0566f
C490 la_data_in[118] la_data_out[118] 0.0566f
C491 wbs_dat_o[28] wbs_adr_i[29] 0.0566f
C492 la_oenb[120] la_data_out[120] 0.0566f
C493 la_oenb[124] la_data_out[124] 0.0566f
C494 io_oeb[8] io_out[8] 0.0824f
C495 io_out[11] a_336716_619863# 0.143f
C496 la_oenb[31] la_data_in[32] 0.0566f
C497 io_oeb[2] io_out[2] 0.0824f
C498 la_data_in[102] la_oenb[101] 0.0566f
C499 la_data_in[22] la_data_out[22] 0.0566f
C500 la_data_out[97] la_oenb[97] 0.0566f
C501 la_oenb[86] la_data_out[86] 0.0566f
C502 io_out[11] gpio_analog[3] 1.33f
C503 a_343294_620745# a_345642_620402# 0.0129f
C504 gpio_noesd[8] io_in_3v3[15] 0.0824f
C505 la_data_out[76] la_oenb[76] 0.0566f
C506 wbs_adr_i[25] wbs_dat_i[25] 0.0566f
C507 la_data_in[14] la_data_out[14] 0.0566f
C508 la_oenb[112] la_data_out[112] 0.0566f
C509 la_data_in[64] la_data_out[64] 0.0566f
C510 la_oenb[122] la_data_in[123] 0.0566f
C511 wbs_adr_i[16] wbs_dat_i[16] 0.0566f
C512 a_345642_617070# pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN 0.00179f
C513 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT 1.47f
C514 a_337674_622496# pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1 0.205f
C515 la_data_out[73] la_data_in[73] 0.0566f
C516 vdda1 a_343294_615747# 1.59f
C517 la_oenb[120] la_data_in[121] 0.0566f
C518 wbs_adr_i[27] wbs_dat_i[27] 0.0566f
C519 io_oeb[25] io_in_3v3[26] 0.0824f
C520 wbs_adr_i[3] wbs_sel_i[2] 0.0566f
C521 la_oenb[121] la_data_in[122] 0.0566f
C522 la_oenb[108] la_data_in[109] 0.0566f
C523 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.493f
C524 la_oenb[104] la_data_in[105] 0.0566f
C525 la_data_out[25] la_data_in[25] 0.0566f
C526 wbs_dat_o[8] wbs_dat_i[8] 0.0566f
C527 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg a_336716_619863# 0.785f
C528 io_out[12] io_oeb[12] 0.0954f
C529 la_data_out[41] la_oenb[41] 0.0566f
C530 wbs_dat_o[12] wbs_adr_i[13] 0.0566f
C531 la_data_out[7] la_data_in[7] 0.0566f
C532 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT w_336471_617254# 0.228f
C533 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN 0.211f
C534 wbs_adr_i[14] wbs_dat_i[14] 0.0566f
C535 wbs_dat_o[20] wbs_adr_i[21] 0.0566f
C536 wbs_dat_i[30] wbs_dat_o[30] 0.0566f
C537 la_oenb[7] la_data_in[8] 0.0566f
C538 io_out[16] io_out[11] 0.0491f
C539 la_data_in[56] la_data_out[56] 0.0566f
C540 la_data_out[68] la_oenb[68] 0.0566f
C541 vccd1 w_336471_617254# 1.82f
C542 la_oenb[80] la_data_out[80] 0.0566f
C543 io_in[19] io_out[19] 0.0824f
C544 la_data_in[63] la_data_out[63] 0.0566f
C545 la_oenb[3] la_data_in[4] 0.0566f
C546 wbs_dat_o[18] wbs_adr_i[19] 0.0566f
C547 wbs_dat_i[25] wbs_dat_o[25] 0.0566f
C548 la_oenb[72] la_data_in[73] 0.0566f
C549 la_data_out[47] la_oenb[47] 0.0566f
C550 io_in[8] io_in_3v3[8] 0.0824f
C551 la_oenb[102] la_data_in[103] 0.0566f
C552 vdda1 gpio_analog[3] 6.98f
C553 wbs_dat_i[26] wbs_dat_o[26] 0.0566f
C554 la_oenb[122] la_data_out[122] 0.0566f
C555 wbs_adr_i[4] wbs_sel_i[3] 0.0566f
C556 wbs_adr_i[2] wbs_sel_i[1] 0.0566f
C557 la_data_in[38] la_data_out[38] 0.0566f
C558 la_oenb[14] la_data_out[14] 0.0566f
C559 la_oenb[32] la_data_in[33] 0.0566f
C560 la_data_out[36] la_oenb[36] 0.0566f
C561 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT vdda1 4.62f
C562 la_data_in[96] la_data_out[96] 0.0566f
C563 la_oenb[10] la_data_in[11] 0.0566f
C564 la_oenb[52] la_data_out[52] 0.0566f
C565 wbs_dat_o[2] wbs_sel_i[2] 0.0566f
C566 la_oenb[79] la_data_in[80] 0.0566f
C567 gpio_noesd[10] io_in_3v3[17] 0.0824f
C568 la_data_out[123] la_data_in[123] 0.0566f
C569 la_oenb[109] la_data_in[110] 0.0566f
C570 wbs_adr_i[1] wbs_sel_i[0] 0.0566f
C571 la_oenb[92] la_data_in[93] 0.0566f
C572 gpio_noesd[5] gpio_analog[5] 0.0824f
C573 la_oenb[43] la_data_in[44] 0.0566f
C574 io_in_3v3[16] io_in[16] 0.0824f
C575 io_oeb[25] io_out[25] 0.0824f
C576 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT 0.00286f
C577 a_337674_622496# pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.00404f
C578 la_data_out[71] la_oenb[71] 0.0566f
C579 gpio_noesd[14] io_in_3v3[21] 0.0824f
C580 io_in_3v3[21] io_in[21] 0.0824f
C581 la_oenb[56] la_data_out[56] 0.0566f
C582 vccd1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1 6.04f
C583 la_data_in[122] la_data_out[122] 0.0566f
C584 la_data_out[15] la_data_in[15] 0.0566f
C585 io_oeb[15] io_out[15] 0.0939f
C586 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT gpio_analog[3] 0.0153f
C587 la_data_in[51] la_data_out[51] 0.0566f
C588 la_oenb[21] la_data_in[22] 0.0566f
C589 la_oenb[50] la_data_out[50] 0.0566f
C590 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN 0.015f
C591 la_data_out[75] la_oenb[75] 0.0566f
C592 la_data_out[7] la_oenb[7] 0.0566f
C593 io_in[25] io_in_3v3[25] 0.0824f
C594 la_oenb[80] la_data_in[81] 0.0566f
C595 la_oenb[84] la_data_in[85] 0.0566f
C596 la_data_in[30] la_data_out[30] 0.0566f
C597 la_data_out[81] la_oenb[81] 0.0566f
C598 la_oenb[33] la_data_in[34] 0.0566f
C599 la_oenb[77] la_data_in[78] 0.0566f
C600 la_data_out[34] la_oenb[34] 0.0566f
C601 la_data_in[74] la_data_out[74] 0.0566f
C602 la_data_in[10] la_data_out[10] 0.0566f
C603 la_data_in[32] la_data_out[32] 0.0566f
C604 la_data_in[106] la_data_out[106] 0.0566f
C605 io_in_3v3[0] io_in[0] 0.0824f
C606 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN 0.105f
C607 wb_rst_i wbs_ack_o 0.0566f
C608 la_data_in[5] la_data_out[5] 0.0566f
C609 la_data_in[92] la_oenb[91] 0.0566f
C610 la_data_out[19] la_oenb[19] 0.0566f
C611 io_out[16] io_oeb[16] 0.095f
C612 la_oenb[96] la_data_in[97] 0.0566f
C613 wbs_dat_i[3] wbs_dat_o[3] 0.0566f
C614 la_oenb[64] la_data_out[64] 0.0566f
C615 gpio_analog[7] gpio_noesd[7] 0.0824f
C616 wbs_dat_i[21] wbs_dat_o[21] 0.0566f
C617 la_oenb[19] la_data_in[20] 0.0566f
C618 la_data_out[123] la_oenb[123] 0.0566f
C619 la_data_in[68] la_oenb[67] 0.0566f
C620 io_in[3] io_in_3v3[3] 0.0824f
C621 la_data_out[99] la_data_in[99] 0.0566f
C622 la_oenb[88] la_data_in[89] 0.0566f
C623 wbs_dat_i[2] wbs_dat_o[2] 0.0566f
C624 io_out[22] io_in[22] 0.0824f
C625 la_data_in[60] la_data_out[60] 0.0566f
C626 la_data_in[20] la_data_out[20] 0.0566f
C627 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN 0.109f
C628 io_oeb[0] io_out[0] 0.0824f
C629 la_data_in[24] la_data_out[24] 0.0566f
C630 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT io_out[12] 0.00182f
C631 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.0712f
C632 a_343294_619079# pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT 0.00155f
C633 la_data_in[27] la_data_out[27] 0.0566f
C634 la_oenb[62] la_data_in[63] 0.0566f
C635 la_oenb[100] la_data_in[101] 0.0566f
C636 a_337674_622496# vccd1 0.511f
C637 vccd1 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT 0.136f
C638 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN a_343294_620745# 0.664f
C639 wbs_dat_o[19] wbs_adr_i[20] 0.0566f
C640 vccd1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 12.6f
C641 la_data_out[30] la_oenb[30] 0.0566f
C642 a_345642_618736# pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT 3.31e-19
C643 la_data_in[11] la_data_out[11] 0.0566f
C644 la_data_out[41] la_data_in[41] 0.0566f
C645 la_oenb[98] la_data_in[99] 0.0566f
C646 io_analog[4] m3_324294_701080# 0.0136f
C647 la_data_in[50] la_data_out[50] 0.0566f
C648 la_data_in[60] la_oenb[59] 0.0566f
C649 io_clamp_high[1] io_analog[5] 0.972f
C650 la_data_out[55] la_oenb[55] 0.0566f
C651 la_oenb[4] la_data_in[5] 0.0566f
C652 la_data_out[25] la_oenb[25] 0.0566f
C653 la_data_out[23] la_oenb[23] 0.0566f
C654 wbs_adr_i[10] wbs_dat_i[10] 0.0566f
C655 io_in_3v3[13] gpio_noesd[6] 0.0824f
C656 io_out[12] io_in[12] 0.0824f
C657 gpio_analog[7] vccd1 2.33f
C658 la_data_in[114] la_data_out[114] 0.0566f
C659 io_out[13] io_in[13] 0.0824f
C660 wbs_adr_i[30] wbs_dat_i[30] 0.0566f
C661 a_343294_620745# vdda1 1.59f
C662 la_data_out[21] la_oenb[21] 0.0566f
C663 la_oenb[95] la_data_in[96] 0.0566f
C664 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN io_out[12] 4.67e-20
C665 gpio_noesd[15] io_in_3v3[22] 0.0824f
C666 la_oenb[24] la_data_in[25] 0.0566f
C667 gpio_analog[14] gpio_noesd[14] 0.0824f
C668 io_out[16] io_out[15] 20.9f
C669 la_data_out[74] la_oenb[74] 0.0566f
C670 la_data_in[4] la_data_out[4] 0.0566f
C671 wbs_dat_o[0] wbs_sel_i[0] 0.0566f
C672 gpio_noesd[0] gpio_analog[0] 0.0824f
C673 wbs_adr_i[2] wbs_dat_i[2] 0.0566f
C674 la_data_out[59] la_oenb[59] 0.0566f
C675 wbs_adr_i[0] wbs_dat_i[0] 0.0566f
C676 gpio_analog[9] gpio_noesd[9] 0.0824f
C677 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN 1.47f
C678 la_data_out[35] la_oenb[35] 0.0566f
C679 la_data_out[31] la_data_in[31] 0.0566f
C680 la_oenb[70] la_data_in[71] 0.0566f
C681 io_out[0] io_in[0] 0.0824f
C682 vccd1 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT 0.328f
C683 io_in[14] io_in_3v3[14] 0.0824f
C684 wbs_dat_i[9] wbs_dat_o[9] 0.0566f
C685 io_in_3v3[17] io_in[17] 0.0824f
C686 io_in_3v3[12] gpio_noesd[5] 0.0824f
C687 la_oenb[18] la_data_out[18] 0.0566f
C688 la_data_out[29] la_oenb[29] 0.0566f
C689 la_data_in[102] la_data_out[102] 0.0566f
C690 la_data_out[113] la_oenb[113] 0.0566f
C691 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN vdda1 4.55f
C692 io_in_3v3[24] gpio_noesd[17] 0.0824f
C693 io_out[12] io_out[11] 28.8f
C694 la_data_out[93] la_oenb[93] 0.0566f
C695 la_data_in[62] la_data_out[62] 0.0566f
C696 io_out[23] io_in[23] 0.0824f
C697 a_343294_620745# pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT 1.07f
C698 la_data_in[126] la_data_out[126] 0.0566f
C699 wbs_dat_o[26] wbs_adr_i[27] 0.0566f
C700 la_oenb[111] la_data_in[112] 0.0566f
C701 la_data_out[116] la_oenb[116] 0.0566f
C702 vdda1 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN 4.57f
C703 io_analog[6] io_clamp_low[2] 0.972f
C704 io_in[25] io_out[25] 0.0824f
C705 la_data_out[109] la_data_in[109] 0.0566f
C706 io_out[14] io_oeb[14] 0.0824f
C707 io_in_3v3[24] io_in[24] 0.0824f
C708 la_data_out[55] la_data_in[55] 0.0566f
C709 gpio_analog[8] gpio_noesd[8] 0.0824f
C710 user_clock2 user_irq[0] 0.0566f
C711 la_oenb[32] la_data_out[32] 0.0566f
C712 la_data_out[69] la_oenb[69] 0.0566f
C713 wbs_adr_i[19] wbs_dat_i[19] 0.0566f
C714 la_data_out[10] la_oenb[10] 0.0566f
C715 la_oenb[117] la_data_in[118] 0.0566f
C716 io_out[2] io_in[2] 0.0824f
C717 a_345642_618736# pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN 1.06e-19
C718 la_data_out[63] la_oenb[63] 0.0566f
C719 io_oeb[9] io_out[9] 0.0824f
C720 vccd1 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT 0.199f
C721 io_out[10] io_oeb[10] 0.0824f
C722 la_data_out[59] la_data_in[59] 0.0566f
C723 la_oenb[48] la_data_in[49] 0.0566f
C724 la_data_out[49] la_data_in[49] 0.0566f
C725 la_data_in[33] la_data_out[33] 0.0566f
C726 io_in_3v3[23] io_in[23] 0.0824f
C727 la_data_out[65] la_oenb[65] 0.0566f
C728 la_data_out[43] la_oenb[43] 0.0566f
C729 wbs_dat_i[17] wbs_dat_o[17] 0.0566f
C730 la_data_in[94] la_data_out[94] 0.0566f
C731 io_oeb[3] io_out[3] 0.0824f
C732 la_oenb[20] la_data_in[21] 0.0566f
C733 io_out[12] vdda1 5.73f
C734 gpio_analog[16] gpio_noesd[16] 0.0824f
C735 wbs_adr_i[13] wbs_dat_i[13] 0.0566f
C736 la_oenb[45] la_data_in[46] 0.0566f
C737 la_oenb[110] la_data_in[111] 0.0566f
C738 wbs_dat_o[13] wbs_adr_i[14] 0.0566f
C739 la_data_out[48] la_oenb[48] 0.0566f
C740 a_345642_617070# pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT 1.09e-19
C741 la_oenb[8] la_data_in[9] 0.0566f
C742 la_oenb[57] la_data_in[58] 0.0566f
C743 la_oenb[6] la_data_in[7] 0.0566f
C744 la_oenb[36] la_data_in[37] 0.0566f
C745 la_data_out[67] la_oenb[67] 0.0566f
C746 la_oenb[38] la_data_in[39] 0.0566f
C747 io_clamp_low[1] m3_225094_700796# 0.00195f
C748 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 3.73e-20
C749 wbs_dat_o[3] wbs_sel_i[3] 0.0566f
C750 la_oenb[8] la_data_out[8] 0.0566f
C751 a_345642_618736# vdda1 1.59f
C752 la_data_in[18] la_data_out[18] 0.0566f
C753 la_data_in[92] la_data_out[92] 0.0566f
C754 la_oenb[108] la_data_out[108] 0.0566f
C755 la_oenb[87] la_data_in[88] 0.0566f
C756 io_out[21] io_oeb[21] 0.0824f
C757 a_345642_620402# pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT 1.22f
C758 la_data_out[78] la_oenb[78] 0.0566f
C759 la_data_out[73] la_oenb[73] 0.0566f
C760 la_data_out[77] la_oenb[77] 0.0566f
C761 la_data_in[106] la_oenb[105] 0.0566f
C762 la_data_in[100] la_data_out[100] 0.0566f
C763 wbs_dat_i[23] wbs_adr_i[23] 0.0566f
C764 a_339370_618592# pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.21f
C765 io_oeb[24] io_out[24] 0.0824f
C766 wbs_dat_i[29] wbs_adr_i[29] 0.0566f
C767 la_data_in[113] la_data_out[113] 0.0566f
C768 la_data_out[95] la_oenb[95] 0.0566f
C769 io_in_3v3[2] io_oeb[1] 0.0824f
C770 la_data_out[66] la_oenb[66] 0.0566f
C771 wbs_adr_i[28] wbs_dat_o[27] 0.0566f
C772 io_out[11] w_336471_617254# 0.219f
C773 a_345642_617070# a_343294_617413# 0.0129f
C774 io_oeb[3] io_in_3v3[4] 0.0824f
C775 a_343294_617413# pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT 1.5e-19
C776 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN a_343294_615747# 1.07f
C777 gpio_analog[3] gpio_noesd[3] 0.0824f
C778 la_oenb[65] la_data_in[66] 0.0566f
C779 la_data_out[58] la_oenb[58] 0.0566f
C780 la_data_out[69] la_data_in[69] 0.0566f
C781 la_data_out[119] la_oenb[119] 0.0566f
C782 la_data_in[70] la_data_out[70] 0.0566f
C783 la_data_in[39] la_data_out[39] 0.0566f
C784 la_data_out[92] la_oenb[92] 0.0566f
C785 wbs_dat_o[14] wbs_adr_i[15] 0.0566f
C786 a_345642_615404# pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT 3.31e-19
C787 la_data_in[84] la_data_out[84] 0.0566f
C788 la_data_out[114] la_oenb[114] 0.0566f
C789 wbs_dat_i[9] wbs_adr_i[9] 0.0566f
C790 la_oenb[13] la_data_in[14] 0.0566f
C791 io_in[20] io_out[20] 0.0824f
C792 la_data_out[4] la_oenb[4] 0.0566f
C793 la_oenb[35] la_data_in[36] 0.0566f
C794 vccd1 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT 0.113f
C795 io_in_3v3[20] io_in[20] 0.0824f
C796 la_oenb[62] la_data_out[62] 0.0566f
C797 io_analog[6] io_clamp_high[2] 0.972f
C798 la_data_in[72] la_oenb[71] 0.0566f
C799 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT 0.113f
C800 a_337674_621712# pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1 0.491f
C801 la_oenb[51] la_data_in[52] 0.0566f
C802 wbs_dat_i[4] wbs_dat_o[4] 0.0566f
C803 la_oenb[20] la_data_out[20] 0.0566f
C804 io_in_3v3[1] io_in[1] 0.0824f
C805 la_oenb[99] la_data_in[100] 0.0566f
C806 m3_170894_700738# io_clamp_high[2] 3.89e-19
C807 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN 0.191f
C808 la_oenb[22] la_data_out[22] 0.0566f
C809 la_oenb[78] la_data_in[79] 0.0566f
C810 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1 io_out[11] 0.00398f
C811 vccd1 a_339370_618592# 0.51f
C812 m3_676_419176# io_out[16] 0.00399f
C813 la_oenb[84] la_data_out[84] 0.0566f
C814 io_analog[4] vssa1 0.324p
C815 io_analog[5] vssa1 23.6f
C816 io_analog[6] vssa1 23.6f
C817 io_in_3v3[0] vssa1 0.507f
C818 io_oeb[26] vssa1 0.507f
C819 io_in[0] vssa1 0.399f
C820 io_out[26] vssa1 0.399f
C821 io_out[0] vssa1 0.399f
C822 io_in[26] vssa1 0.399f
C823 io_oeb[0] vssa1 0.399f
C824 io_in_3v3[26] vssa1 0.399f
C825 io_in_3v3[1] vssa1 0.399f
C826 io_oeb[25] vssa1 0.399f
C827 io_in[1] vssa1 0.399f
C828 io_out[25] vssa1 0.399f
C829 io_out[1] vssa1 0.399f
C830 io_in[25] vssa1 0.399f
C831 io_oeb[1] vssa1 0.399f
C832 io_in_3v3[25] vssa1 0.399f
C833 io_in_3v3[2] vssa1 0.399f
C834 io_oeb[24] vssa1 0.399f
C835 io_in[2] vssa1 0.399f
C836 io_out[24] vssa1 0.399f
C837 io_out[2] vssa1 0.399f
C838 io_in[24] vssa1 0.399f
C839 io_oeb[2] vssa1 0.399f
C840 io_in_3v3[24] vssa1 0.399f
C841 io_in_3v3[3] vssa1 0.399f
C842 gpio_noesd[17] vssa1 0.399f
C843 io_in[3] vssa1 0.399f
C844 gpio_analog[17] vssa1 0.507f
C845 io_out[3] vssa1 0.399f
C846 io_oeb[3] vssa1 0.399f
C847 io_in_3v3[4] vssa1 0.399f
C848 io_in[4] vssa1 0.399f
C849 io_out[4] vssa1 0.399f
C850 io_oeb[4] vssa1 0.507f
C851 io_oeb[23] vssa1 0.507f
C852 io_out[23] vssa1 0.399f
C853 io_in[23] vssa1 0.399f
C854 io_in_3v3[23] vssa1 0.399f
C855 gpio_noesd[16] vssa1 0.399f
C856 gpio_analog[16] vssa1 0.507f
C857 io_in_3v3[5] vssa1 0.507f
C858 io_in[5] vssa1 0.399f
C859 io_out[5] vssa1 0.399f
C860 io_oeb[5] vssa1 0.507f
C861 io_oeb[22] vssa1 0.507f
C862 io_out[22] vssa1 0.399f
C863 io_in[22] vssa1 0.399f
C864 io_in_3v3[22] vssa1 0.399f
C865 gpio_noesd[15] vssa1 0.399f
C866 gpio_analog[15] vssa1 0.507f
C867 io_in_3v3[6] vssa1 0.507f
C868 io_in[6] vssa1 0.399f
C869 io_out[6] vssa1 0.399f
C870 io_oeb[6] vssa1 0.507f
C871 io_oeb[21] vssa1 0.507f
C872 io_out[21] vssa1 0.399f
C873 io_in[21] vssa1 0.399f
C874 io_in_3v3[21] vssa1 0.399f
C875 gpio_noesd[14] vssa1 0.399f
C876 gpio_analog[14] vssa1 0.507f
C877 vssd2 vssa1 13.3f
C878 vdda2 vssa1 13.3f
C879 io_oeb[20] vssa1 0.507f
C880 io_out[20] vssa1 0.399f
C881 io_in[20] vssa1 0.399f
C882 io_in_3v3[20] vssa1 0.399f
C883 gpio_noesd[13] vssa1 0.399f
C884 gpio_analog[13] vssa1 0.507f
C885 gpio_analog[0] vssa1 0.507f
C886 gpio_noesd[0] vssa1 0.399f
C887 io_in_3v3[7] vssa1 0.399f
C888 io_in[7] vssa1 0.399f
C889 io_out[7] vssa1 0.399f
C890 io_oeb[7] vssa1 0.507f
C891 io_oeb[19] vssa1 0.507f
C892 io_out[19] vssa1 0.399f
C893 io_in[19] vssa1 0.399f
C894 io_in_3v3[19] vssa1 0.399f
C895 gpio_noesd[12] vssa1 0.399f
C896 gpio_analog[12] vssa1 0.507f
C897 gpio_analog[1] vssa1 0.507f
C898 gpio_noesd[1] vssa1 0.399f
C899 io_in_3v3[8] vssa1 0.399f
C900 io_in[8] vssa1 0.399f
C901 io_out[8] vssa1 0.399f
C902 io_oeb[8] vssa1 0.507f
C903 io_oeb[18] vssa1 0.507f
C904 io_out[18] vssa1 0.399f
C905 io_in[18] vssa1 0.399f
C906 io_in_3v3[18] vssa1 0.399f
C907 gpio_noesd[11] vssa1 0.399f
C908 gpio_analog[11] vssa1 0.507f
C909 gpio_analog[2] vssa1 0.507f
C910 gpio_noesd[2] vssa1 0.399f
C911 io_in_3v3[9] vssa1 0.399f
C912 io_in[9] vssa1 0.399f
C913 io_out[9] vssa1 0.399f
C914 io_oeb[9] vssa1 0.507f
C915 io_oeb[17] vssa1 0.507f
C916 io_out[17] vssa1 0.399f
C917 io_in[17] vssa1 0.399f
C918 io_in_3v3[17] vssa1 0.399f
C919 gpio_noesd[10] vssa1 0.399f
C920 gpio_analog[10] vssa1 0.507f
C921 gpio_noesd[3] vssa1 0.399f
C922 io_in_3v3[10] vssa1 0.399f
C923 io_in[10] vssa1 0.399f
C924 io_out[10] vssa1 0.399f
C925 io_oeb[10] vssa1 0.507f
C926 gpio_analog[4] vssa1 0.507f
C927 gpio_noesd[4] vssa1 0.399f
C928 io_in_3v3[11] vssa1 0.399f
C929 io_in[11] vssa1 0.399f
C930 io_oeb[11] vssa1 0.565f
C931 gpio_analog[5] vssa1 0.507f
C932 gpio_noesd[5] vssa1 0.399f
C933 io_in_3v3[12] vssa1 0.399f
C934 io_in[12] vssa1 0.399f
C935 io_oeb[12] vssa1 0.557f
C936 gpio_analog[6] vssa1 0.507f
C937 gpio_noesd[6] vssa1 0.399f
C938 io_in_3v3[13] vssa1 0.399f
C939 io_in[13] vssa1 0.399f
C940 io_out[13] vssa1 0.399f
C941 io_oeb[13] vssa1 0.507f
C942 io_oeb[16] vssa1 0.554f
C943 io_in[16] vssa1 0.399f
C944 io_in_3v3[16] vssa1 0.399f
C945 gpio_noesd[9] vssa1 0.399f
C946 gpio_analog[9] vssa1 0.507f
C947 io_oeb[15] vssa1 0.549f
C948 io_in[15] vssa1 0.399f
C949 io_in_3v3[15] vssa1 0.399f
C950 gpio_noesd[8] vssa1 0.399f
C951 gpio_analog[8] vssa1 0.507f
C952 io_oeb[14] vssa1 0.507f
C953 io_out[14] vssa1 0.399f
C954 io_in[14] vssa1 0.399f
C955 io_in_3v3[14] vssa1 0.399f
C956 gpio_noesd[7] vssa1 0.399f
C957 vssa2 vssa1 13.3f
C958 vccd2 vssa1 13.3f
C959 io_analog[0] vssa1 6.94f
C960 io_analog[1] vssa1 6.94f
C961 io_analog[2] vssa1 6.94f
C962 io_analog[3] vssa1 6.94f
C963 io_clamp_high[0] vssa1 3.27f
C964 io_clamp_low[0] vssa1 3.29f
C965 io_clamp_high[1] vssa1 3.74f
C966 io_clamp_low[1] vssa1 3.75f
C967 io_clamp_high[2] vssa1 3.79f
C968 io_analog[10] vssa1 6.94f
C969 io_clamp_low[2] vssa1 3.79f
C970 io_analog[7] vssa1 6.94f
C971 io_analog[8] vssa1 6.94f
C972 io_analog[9] vssa1 6.94f
C973 user_irq[2] vssa1 0.513f
C974 user_irq[1] vssa1 0.437f
C975 user_irq[0] vssa1 0.437f
C976 user_clock2 vssa1 0.437f
C977 la_oenb[127] vssa1 0.437f
C978 la_data_out[127] vssa1 0.437f
C979 la_data_in[127] vssa1 0.437f
C980 la_oenb[126] vssa1 0.437f
C981 la_data_out[126] vssa1 0.437f
C982 la_data_in[126] vssa1 0.437f
C983 la_oenb[125] vssa1 0.437f
C984 la_data_out[125] vssa1 0.437f
C985 la_data_in[125] vssa1 0.437f
C986 la_oenb[124] vssa1 0.437f
C987 la_data_out[124] vssa1 0.437f
C988 la_data_in[124] vssa1 0.437f
C989 la_oenb[123] vssa1 0.437f
C990 la_data_out[123] vssa1 0.437f
C991 la_data_in[123] vssa1 0.437f
C992 la_oenb[122] vssa1 0.437f
C993 la_data_out[122] vssa1 0.437f
C994 la_data_in[122] vssa1 0.437f
C995 la_oenb[121] vssa1 0.437f
C996 la_data_out[121] vssa1 0.437f
C997 la_data_in[121] vssa1 0.437f
C998 la_oenb[120] vssa1 0.437f
C999 la_data_out[120] vssa1 0.437f
C1000 la_data_in[120] vssa1 0.437f
C1001 la_oenb[119] vssa1 0.437f
C1002 la_data_out[119] vssa1 0.437f
C1003 la_data_in[119] vssa1 0.437f
C1004 la_oenb[118] vssa1 0.437f
C1005 la_data_out[118] vssa1 0.437f
C1006 la_data_in[118] vssa1 0.437f
C1007 la_oenb[117] vssa1 0.437f
C1008 la_data_out[117] vssa1 0.437f
C1009 la_data_in[117] vssa1 0.437f
C1010 la_oenb[116] vssa1 0.437f
C1011 la_data_out[116] vssa1 0.437f
C1012 la_data_in[116] vssa1 0.437f
C1013 la_oenb[115] vssa1 0.437f
C1014 la_data_out[115] vssa1 0.437f
C1015 la_data_in[115] vssa1 0.437f
C1016 la_oenb[114] vssa1 0.437f
C1017 la_data_out[114] vssa1 0.437f
C1018 la_data_in[114] vssa1 0.437f
C1019 la_oenb[113] vssa1 0.437f
C1020 la_data_out[113] vssa1 0.437f
C1021 la_data_in[113] vssa1 0.437f
C1022 la_oenb[112] vssa1 0.437f
C1023 la_data_out[112] vssa1 0.437f
C1024 la_data_in[112] vssa1 0.437f
C1025 la_oenb[111] vssa1 0.437f
C1026 la_data_out[111] vssa1 0.437f
C1027 la_data_in[111] vssa1 0.437f
C1028 la_oenb[110] vssa1 0.437f
C1029 la_data_out[110] vssa1 0.437f
C1030 la_data_in[110] vssa1 0.437f
C1031 la_oenb[109] vssa1 0.437f
C1032 la_data_out[109] vssa1 0.437f
C1033 la_data_in[109] vssa1 0.437f
C1034 la_oenb[108] vssa1 0.437f
C1035 la_data_out[108] vssa1 0.437f
C1036 la_data_in[108] vssa1 0.437f
C1037 la_oenb[107] vssa1 0.437f
C1038 la_data_out[107] vssa1 0.437f
C1039 la_data_in[107] vssa1 0.437f
C1040 la_oenb[106] vssa1 0.437f
C1041 la_data_out[106] vssa1 0.437f
C1042 la_data_in[106] vssa1 0.437f
C1043 la_oenb[105] vssa1 0.437f
C1044 la_data_out[105] vssa1 0.437f
C1045 la_data_in[105] vssa1 0.437f
C1046 la_oenb[104] vssa1 0.437f
C1047 la_data_out[104] vssa1 0.437f
C1048 la_data_in[104] vssa1 0.437f
C1049 la_oenb[103] vssa1 0.437f
C1050 la_data_out[103] vssa1 0.437f
C1051 la_data_in[103] vssa1 0.437f
C1052 la_oenb[102] vssa1 0.437f
C1053 la_data_out[102] vssa1 0.437f
C1054 la_data_in[102] vssa1 0.437f
C1055 la_oenb[101] vssa1 0.437f
C1056 la_data_out[101] vssa1 0.437f
C1057 la_data_in[101] vssa1 0.437f
C1058 la_oenb[100] vssa1 0.437f
C1059 la_data_out[100] vssa1 0.437f
C1060 la_data_in[100] vssa1 0.437f
C1061 la_oenb[99] vssa1 0.437f
C1062 la_data_out[99] vssa1 0.437f
C1063 la_data_in[99] vssa1 0.437f
C1064 la_oenb[98] vssa1 0.437f
C1065 la_data_out[98] vssa1 0.437f
C1066 la_data_in[98] vssa1 0.437f
C1067 la_oenb[97] vssa1 0.437f
C1068 la_data_out[97] vssa1 0.437f
C1069 la_data_in[97] vssa1 0.437f
C1070 la_oenb[96] vssa1 0.437f
C1071 la_data_out[96] vssa1 0.437f
C1072 la_data_in[96] vssa1 0.437f
C1073 la_oenb[95] vssa1 0.437f
C1074 la_data_out[95] vssa1 0.437f
C1075 la_data_in[95] vssa1 0.437f
C1076 la_oenb[94] vssa1 0.437f
C1077 la_data_out[94] vssa1 0.437f
C1078 la_data_in[94] vssa1 0.437f
C1079 la_oenb[93] vssa1 0.437f
C1080 la_data_out[93] vssa1 0.437f
C1081 la_data_in[93] vssa1 0.437f
C1082 la_oenb[92] vssa1 0.437f
C1083 la_data_out[92] vssa1 0.437f
C1084 la_data_in[92] vssa1 0.437f
C1085 la_oenb[91] vssa1 0.437f
C1086 la_data_out[91] vssa1 0.437f
C1087 la_data_in[91] vssa1 0.437f
C1088 la_oenb[90] vssa1 0.437f
C1089 la_data_out[90] vssa1 0.437f
C1090 la_data_in[90] vssa1 0.437f
C1091 la_oenb[89] vssa1 0.437f
C1092 la_data_out[89] vssa1 0.437f
C1093 la_data_in[89] vssa1 0.437f
C1094 la_oenb[88] vssa1 0.437f
C1095 la_data_out[88] vssa1 0.437f
C1096 la_data_in[88] vssa1 0.437f
C1097 la_oenb[87] vssa1 0.437f
C1098 la_data_out[87] vssa1 0.437f
C1099 la_data_in[87] vssa1 0.437f
C1100 la_oenb[86] vssa1 0.437f
C1101 la_data_out[86] vssa1 0.437f
C1102 la_data_in[86] vssa1 0.437f
C1103 la_oenb[85] vssa1 0.437f
C1104 la_data_out[85] vssa1 0.437f
C1105 la_data_in[85] vssa1 0.437f
C1106 la_oenb[84] vssa1 0.437f
C1107 la_data_out[84] vssa1 0.437f
C1108 la_data_in[84] vssa1 0.437f
C1109 la_oenb[83] vssa1 0.437f
C1110 la_data_out[83] vssa1 0.437f
C1111 la_data_in[83] vssa1 0.437f
C1112 la_oenb[82] vssa1 0.437f
C1113 la_data_out[82] vssa1 0.437f
C1114 la_data_in[82] vssa1 0.437f
C1115 la_oenb[81] vssa1 0.437f
C1116 la_data_out[81] vssa1 0.437f
C1117 la_data_in[81] vssa1 0.437f
C1118 la_oenb[80] vssa1 0.437f
C1119 la_data_out[80] vssa1 0.437f
C1120 la_data_in[80] vssa1 0.437f
C1121 la_oenb[79] vssa1 0.437f
C1122 la_data_out[79] vssa1 0.437f
C1123 la_data_in[79] vssa1 0.437f
C1124 la_oenb[78] vssa1 0.437f
C1125 la_data_out[78] vssa1 0.437f
C1126 la_data_in[78] vssa1 0.437f
C1127 la_oenb[77] vssa1 0.437f
C1128 la_data_out[77] vssa1 0.437f
C1129 la_data_in[77] vssa1 0.437f
C1130 la_oenb[76] vssa1 0.437f
C1131 la_data_out[76] vssa1 0.437f
C1132 la_data_in[76] vssa1 0.437f
C1133 la_oenb[75] vssa1 0.437f
C1134 la_data_out[75] vssa1 0.437f
C1135 la_data_in[75] vssa1 0.437f
C1136 la_oenb[74] vssa1 0.437f
C1137 la_data_out[74] vssa1 0.437f
C1138 la_data_in[74] vssa1 0.437f
C1139 la_oenb[73] vssa1 0.437f
C1140 la_data_out[73] vssa1 0.437f
C1141 la_data_in[73] vssa1 0.437f
C1142 la_oenb[72] vssa1 0.437f
C1143 la_data_out[72] vssa1 0.437f
C1144 la_data_in[72] vssa1 0.437f
C1145 la_oenb[71] vssa1 0.437f
C1146 la_data_out[71] vssa1 0.437f
C1147 la_data_in[71] vssa1 0.437f
C1148 la_oenb[70] vssa1 0.437f
C1149 la_data_out[70] vssa1 0.437f
C1150 la_data_in[70] vssa1 0.437f
C1151 la_oenb[69] vssa1 0.437f
C1152 la_data_out[69] vssa1 0.437f
C1153 la_data_in[69] vssa1 0.437f
C1154 la_oenb[68] vssa1 0.437f
C1155 la_data_out[68] vssa1 0.437f
C1156 la_data_in[68] vssa1 0.437f
C1157 la_oenb[67] vssa1 0.437f
C1158 la_data_out[67] vssa1 0.437f
C1159 la_data_in[67] vssa1 0.437f
C1160 la_oenb[66] vssa1 0.437f
C1161 la_data_out[66] vssa1 0.437f
C1162 la_data_in[66] vssa1 0.437f
C1163 la_oenb[65] vssa1 0.437f
C1164 la_data_out[65] vssa1 0.437f
C1165 la_data_in[65] vssa1 0.437f
C1166 la_oenb[64] vssa1 0.437f
C1167 la_data_out[64] vssa1 0.437f
C1168 la_data_in[64] vssa1 0.437f
C1169 la_oenb[63] vssa1 0.437f
C1170 la_data_out[63] vssa1 0.437f
C1171 la_data_in[63] vssa1 0.437f
C1172 la_oenb[62] vssa1 0.437f
C1173 la_data_out[62] vssa1 0.437f
C1174 la_data_in[62] vssa1 0.437f
C1175 la_oenb[61] vssa1 0.437f
C1176 la_data_out[61] vssa1 0.437f
C1177 la_data_in[61] vssa1 0.437f
C1178 la_oenb[60] vssa1 0.437f
C1179 la_data_out[60] vssa1 0.437f
C1180 la_data_in[60] vssa1 0.437f
C1181 la_oenb[59] vssa1 0.437f
C1182 la_data_out[59] vssa1 0.437f
C1183 la_data_in[59] vssa1 0.437f
C1184 la_oenb[58] vssa1 0.437f
C1185 la_data_out[58] vssa1 0.437f
C1186 la_data_in[58] vssa1 0.437f
C1187 la_oenb[57] vssa1 0.437f
C1188 la_data_out[57] vssa1 0.437f
C1189 la_data_in[57] vssa1 0.437f
C1190 la_oenb[56] vssa1 0.437f
C1191 la_data_out[56] vssa1 0.437f
C1192 la_data_in[56] vssa1 0.437f
C1193 la_oenb[55] vssa1 0.437f
C1194 la_data_out[55] vssa1 0.437f
C1195 la_data_in[55] vssa1 0.437f
C1196 la_oenb[54] vssa1 0.437f
C1197 la_data_out[54] vssa1 0.437f
C1198 la_data_in[54] vssa1 0.437f
C1199 la_oenb[53] vssa1 0.437f
C1200 la_data_out[53] vssa1 0.437f
C1201 la_data_in[53] vssa1 0.437f
C1202 la_oenb[52] vssa1 0.437f
C1203 la_data_out[52] vssa1 0.437f
C1204 la_data_in[52] vssa1 0.437f
C1205 la_oenb[51] vssa1 0.437f
C1206 la_data_out[51] vssa1 0.437f
C1207 la_data_in[51] vssa1 0.437f
C1208 la_oenb[50] vssa1 0.437f
C1209 la_data_out[50] vssa1 0.437f
C1210 la_data_in[50] vssa1 0.437f
C1211 la_oenb[49] vssa1 0.437f
C1212 la_data_out[49] vssa1 0.437f
C1213 la_data_in[49] vssa1 0.437f
C1214 la_oenb[48] vssa1 0.437f
C1215 la_data_out[48] vssa1 0.437f
C1216 la_data_in[48] vssa1 0.437f
C1217 la_oenb[47] vssa1 0.437f
C1218 la_data_out[47] vssa1 0.437f
C1219 la_data_in[47] vssa1 0.437f
C1220 la_oenb[46] vssa1 0.437f
C1221 la_data_out[46] vssa1 0.437f
C1222 la_data_in[46] vssa1 0.437f
C1223 la_oenb[45] vssa1 0.437f
C1224 la_data_out[45] vssa1 0.437f
C1225 la_data_in[45] vssa1 0.437f
C1226 la_oenb[44] vssa1 0.437f
C1227 la_data_out[44] vssa1 0.437f
C1228 la_data_in[44] vssa1 0.437f
C1229 la_oenb[43] vssa1 0.437f
C1230 la_data_out[43] vssa1 0.437f
C1231 la_data_in[43] vssa1 0.437f
C1232 la_oenb[42] vssa1 0.437f
C1233 la_data_out[42] vssa1 0.437f
C1234 la_data_in[42] vssa1 0.437f
C1235 la_oenb[41] vssa1 0.437f
C1236 la_data_out[41] vssa1 0.437f
C1237 la_data_in[41] vssa1 0.437f
C1238 la_oenb[40] vssa1 0.437f
C1239 la_data_out[40] vssa1 0.437f
C1240 la_data_in[40] vssa1 0.437f
C1241 la_oenb[39] vssa1 0.437f
C1242 la_data_out[39] vssa1 0.437f
C1243 la_data_in[39] vssa1 0.437f
C1244 la_oenb[38] vssa1 0.437f
C1245 la_data_out[38] vssa1 0.437f
C1246 la_data_in[38] vssa1 0.437f
C1247 la_oenb[37] vssa1 0.437f
C1248 la_data_out[37] vssa1 0.437f
C1249 la_data_in[37] vssa1 0.437f
C1250 la_oenb[36] vssa1 0.437f
C1251 la_data_out[36] vssa1 0.437f
C1252 la_data_in[36] vssa1 0.437f
C1253 la_oenb[35] vssa1 0.437f
C1254 la_data_out[35] vssa1 0.437f
C1255 la_data_in[35] vssa1 0.437f
C1256 la_oenb[34] vssa1 0.437f
C1257 la_data_out[34] vssa1 0.437f
C1258 la_data_in[34] vssa1 0.437f
C1259 la_oenb[33] vssa1 0.437f
C1260 la_data_out[33] vssa1 0.437f
C1261 la_data_in[33] vssa1 0.437f
C1262 la_oenb[32] vssa1 0.437f
C1263 la_data_out[32] vssa1 0.437f
C1264 la_data_in[32] vssa1 0.437f
C1265 la_oenb[31] vssa1 0.437f
C1266 la_data_out[31] vssa1 0.437f
C1267 la_data_in[31] vssa1 0.437f
C1268 la_oenb[30] vssa1 0.437f
C1269 la_data_out[30] vssa1 0.437f
C1270 la_data_in[30] vssa1 0.437f
C1271 la_oenb[29] vssa1 0.437f
C1272 la_data_out[29] vssa1 0.437f
C1273 la_data_in[29] vssa1 0.437f
C1274 la_oenb[28] vssa1 0.437f
C1275 la_data_out[28] vssa1 0.437f
C1276 la_data_in[28] vssa1 0.437f
C1277 la_oenb[27] vssa1 0.437f
C1278 la_data_out[27] vssa1 0.437f
C1279 la_data_in[27] vssa1 0.437f
C1280 la_oenb[26] vssa1 0.437f
C1281 la_data_out[26] vssa1 0.437f
C1282 la_data_in[26] vssa1 0.437f
C1283 la_oenb[25] vssa1 0.437f
C1284 la_data_out[25] vssa1 0.437f
C1285 la_data_in[25] vssa1 0.437f
C1286 la_oenb[24] vssa1 0.437f
C1287 la_data_out[24] vssa1 0.437f
C1288 la_data_in[24] vssa1 0.437f
C1289 la_oenb[23] vssa1 0.437f
C1290 la_data_out[23] vssa1 0.437f
C1291 la_data_in[23] vssa1 0.437f
C1292 la_oenb[22] vssa1 0.437f
C1293 la_data_out[22] vssa1 0.437f
C1294 la_data_in[22] vssa1 0.437f
C1295 la_oenb[21] vssa1 0.437f
C1296 la_data_out[21] vssa1 0.437f
C1297 la_data_in[21] vssa1 0.437f
C1298 la_oenb[20] vssa1 0.437f
C1299 la_data_out[20] vssa1 0.437f
C1300 la_data_in[20] vssa1 0.437f
C1301 la_oenb[19] vssa1 0.437f
C1302 la_data_out[19] vssa1 0.437f
C1303 la_data_in[19] vssa1 0.437f
C1304 la_oenb[18] vssa1 0.437f
C1305 la_data_out[18] vssa1 0.437f
C1306 la_data_in[18] vssa1 0.437f
C1307 la_oenb[17] vssa1 0.437f
C1308 la_data_out[17] vssa1 0.437f
C1309 la_data_in[17] vssa1 0.437f
C1310 la_oenb[16] vssa1 0.437f
C1311 la_data_out[16] vssa1 0.437f
C1312 la_data_in[16] vssa1 0.437f
C1313 la_oenb[15] vssa1 0.437f
C1314 la_data_out[15] vssa1 0.437f
C1315 la_data_in[15] vssa1 0.437f
C1316 la_oenb[14] vssa1 0.437f
C1317 la_data_out[14] vssa1 0.437f
C1318 la_data_in[14] vssa1 0.437f
C1319 la_oenb[13] vssa1 0.437f
C1320 la_data_out[13] vssa1 0.437f
C1321 la_data_in[13] vssa1 0.437f
C1322 la_oenb[12] vssa1 0.437f
C1323 la_data_out[12] vssa1 0.437f
C1324 la_data_in[12] vssa1 0.437f
C1325 la_oenb[11] vssa1 0.437f
C1326 la_data_out[11] vssa1 0.437f
C1327 la_data_in[11] vssa1 0.437f
C1328 la_oenb[10] vssa1 0.437f
C1329 la_data_out[10] vssa1 0.437f
C1330 la_data_in[10] vssa1 0.437f
C1331 la_oenb[9] vssa1 0.437f
C1332 la_data_out[9] vssa1 0.437f
C1333 la_data_in[9] vssa1 0.437f
C1334 la_oenb[8] vssa1 0.437f
C1335 la_data_out[8] vssa1 0.437f
C1336 la_data_in[8] vssa1 0.437f
C1337 la_oenb[7] vssa1 0.437f
C1338 la_data_out[7] vssa1 0.437f
C1339 la_data_in[7] vssa1 0.437f
C1340 la_oenb[6] vssa1 0.437f
C1341 la_data_out[6] vssa1 0.437f
C1342 la_data_in[6] vssa1 0.437f
C1343 la_oenb[5] vssa1 0.437f
C1344 la_data_out[5] vssa1 0.437f
C1345 la_data_in[5] vssa1 0.437f
C1346 la_oenb[4] vssa1 0.437f
C1347 la_data_out[4] vssa1 0.437f
C1348 la_data_in[4] vssa1 0.437f
C1349 la_oenb[3] vssa1 0.437f
C1350 la_data_out[3] vssa1 0.437f
C1351 la_data_in[3] vssa1 0.437f
C1352 la_oenb[2] vssa1 0.437f
C1353 la_data_out[2] vssa1 0.437f
C1354 la_data_in[2] vssa1 0.437f
C1355 la_oenb[1] vssa1 0.437f
C1356 la_data_out[1] vssa1 0.437f
C1357 la_data_in[1] vssa1 0.437f
C1358 la_oenb[0] vssa1 0.437f
C1359 la_data_out[0] vssa1 0.437f
C1360 la_data_in[0] vssa1 0.437f
C1361 wbs_dat_o[31] vssa1 0.437f
C1362 wbs_dat_i[31] vssa1 0.437f
C1363 wbs_adr_i[31] vssa1 0.437f
C1364 wbs_dat_o[30] vssa1 0.437f
C1365 wbs_dat_i[30] vssa1 0.437f
C1366 wbs_adr_i[30] vssa1 0.437f
C1367 wbs_dat_o[29] vssa1 0.437f
C1368 wbs_dat_i[29] vssa1 0.437f
C1369 wbs_adr_i[29] vssa1 0.437f
C1370 wbs_dat_o[28] vssa1 0.437f
C1371 wbs_dat_i[28] vssa1 0.437f
C1372 wbs_adr_i[28] vssa1 0.437f
C1373 wbs_dat_o[27] vssa1 0.437f
C1374 wbs_dat_i[27] vssa1 0.437f
C1375 wbs_adr_i[27] vssa1 0.437f
C1376 wbs_dat_o[26] vssa1 0.437f
C1377 wbs_dat_i[26] vssa1 0.437f
C1378 wbs_adr_i[26] vssa1 0.437f
C1379 wbs_dat_o[25] vssa1 0.437f
C1380 wbs_dat_i[25] vssa1 0.437f
C1381 wbs_adr_i[25] vssa1 0.437f
C1382 wbs_dat_o[24] vssa1 0.437f
C1383 wbs_dat_i[24] vssa1 0.437f
C1384 wbs_adr_i[24] vssa1 0.437f
C1385 wbs_dat_o[23] vssa1 0.437f
C1386 wbs_dat_i[23] vssa1 0.437f
C1387 wbs_adr_i[23] vssa1 0.437f
C1388 wbs_dat_o[22] vssa1 0.437f
C1389 wbs_dat_i[22] vssa1 0.437f
C1390 wbs_adr_i[22] vssa1 0.437f
C1391 wbs_dat_o[21] vssa1 0.437f
C1392 wbs_dat_i[21] vssa1 0.437f
C1393 wbs_adr_i[21] vssa1 0.437f
C1394 wbs_dat_o[20] vssa1 0.437f
C1395 wbs_dat_i[20] vssa1 0.437f
C1396 wbs_adr_i[20] vssa1 0.437f
C1397 wbs_dat_o[19] vssa1 0.437f
C1398 wbs_dat_i[19] vssa1 0.437f
C1399 wbs_adr_i[19] vssa1 0.437f
C1400 wbs_dat_o[18] vssa1 0.437f
C1401 wbs_dat_i[18] vssa1 0.437f
C1402 wbs_adr_i[18] vssa1 0.437f
C1403 wbs_dat_o[17] vssa1 0.437f
C1404 wbs_dat_i[17] vssa1 0.437f
C1405 wbs_adr_i[17] vssa1 0.437f
C1406 wbs_dat_o[16] vssa1 0.437f
C1407 wbs_dat_i[16] vssa1 0.437f
C1408 wbs_adr_i[16] vssa1 0.437f
C1409 wbs_dat_o[15] vssa1 0.437f
C1410 wbs_dat_i[15] vssa1 0.437f
C1411 wbs_adr_i[15] vssa1 0.437f
C1412 wbs_dat_o[14] vssa1 0.437f
C1413 wbs_dat_i[14] vssa1 0.437f
C1414 wbs_adr_i[14] vssa1 0.437f
C1415 wbs_dat_o[13] vssa1 0.437f
C1416 wbs_dat_i[13] vssa1 0.437f
C1417 wbs_adr_i[13] vssa1 0.437f
C1418 wbs_dat_o[12] vssa1 0.437f
C1419 wbs_dat_i[12] vssa1 0.437f
C1420 wbs_adr_i[12] vssa1 0.437f
C1421 wbs_dat_o[11] vssa1 0.437f
C1422 wbs_dat_i[11] vssa1 0.437f
C1423 wbs_adr_i[11] vssa1 0.437f
C1424 wbs_dat_o[10] vssa1 0.437f
C1425 wbs_dat_i[10] vssa1 0.437f
C1426 wbs_adr_i[10] vssa1 0.437f
C1427 wbs_dat_o[9] vssa1 0.437f
C1428 wbs_dat_i[9] vssa1 0.437f
C1429 wbs_adr_i[9] vssa1 0.437f
C1430 wbs_dat_o[8] vssa1 0.437f
C1431 wbs_dat_i[8] vssa1 0.437f
C1432 wbs_adr_i[8] vssa1 0.437f
C1433 wbs_dat_o[7] vssa1 0.437f
C1434 wbs_dat_i[7] vssa1 0.437f
C1435 wbs_adr_i[7] vssa1 0.437f
C1436 wbs_dat_o[6] vssa1 0.437f
C1437 wbs_dat_i[6] vssa1 0.437f
C1438 wbs_adr_i[6] vssa1 0.437f
C1439 wbs_dat_o[5] vssa1 0.437f
C1440 wbs_dat_i[5] vssa1 0.437f
C1441 wbs_adr_i[5] vssa1 0.437f
C1442 wbs_dat_o[4] vssa1 0.437f
C1443 wbs_dat_i[4] vssa1 0.437f
C1444 wbs_adr_i[4] vssa1 0.437f
C1445 wbs_sel_i[3] vssa1 0.437f
C1446 wbs_dat_o[3] vssa1 0.437f
C1447 wbs_dat_i[3] vssa1 0.437f
C1448 wbs_adr_i[3] vssa1 0.437f
C1449 wbs_sel_i[2] vssa1 0.437f
C1450 wbs_dat_o[2] vssa1 0.437f
C1451 wbs_dat_i[2] vssa1 0.437f
C1452 wbs_adr_i[2] vssa1 0.437f
C1453 wbs_sel_i[1] vssa1 0.437f
C1454 wbs_dat_o[1] vssa1 0.437f
C1455 wbs_dat_i[1] vssa1 0.437f
C1456 wbs_adr_i[1] vssa1 0.437f
C1457 wbs_sel_i[0] vssa1 0.437f
C1458 wbs_dat_o[0] vssa1 0.437f
C1459 wbs_dat_i[0] vssa1 0.437f
C1460 wbs_adr_i[0] vssa1 0.437f
C1461 wbs_we_i vssa1 0.437f
C1462 wbs_stb_i vssa1 0.437f
C1463 wbs_cyc_i vssa1 0.437f
C1464 wbs_ack_o vssa1 0.437f
C1465 wb_rst_i vssa1 0.437f
C1466 wb_clk_i vssa1 0.513f
C1467 m3_583180_455628# vssa1 0.0418f $ **FLOATING
C1468 m3_583220_500050# vssa1 0.0353f $ **FLOATING
C1469 m3_676_419176# vssa1 0.0223f $ **FLOATING
C1470 vssd1 vssa1 1.77p
C1471 m3_660_462398# vssa1 0.0432f $ **FLOATING
C1472 m3_326794_701100# vssa1 0.0387f $ **FLOATING
C1473 m3_324294_701080# vssa1 0.0387f $ **FLOATING
C1474 m3_225094_700796# vssa1 0.0466f $ **FLOATING
C1475 m3_222594_700786# vssa1 0.0485f $ **FLOATING
C1476 m3_173394_700736# vssa1 0.047f $ **FLOATING
C1477 m3_170894_700738# vssa1 0.0466f $ **FLOATING
C1478 gpio_analog[7] vssa1 0.208p
C1479 io_out[16] vssa1 0.242p
C1480 io_out[12] vssa1 0.153p
C1481 a_345642_613738# vssa1 0.41f
C1482 a_343294_614081# vssa1 0.41f
C1483 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT vssa1 8.68f
C1484 a_345642_615404# vssa1 0.41f
C1485 pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN vssa1 8.18f
C1486 a_343294_615747# vssa1 0.41f
C1487 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT vssa1 8.17f
C1488 a_345642_617070# vssa1 0.41f
C1489 pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT vssa1 8.13f
C1490 a_343294_617413# vssa1 0.41f
C1491 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN vssa1 8.5f
C1492 a_345642_618736# vssa1 0.41f
C1493 pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT vssa1 8.14f
C1494 a_343294_619079# vssa1 0.41f
C1495 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN vssa1 8.22f
C1496 a_345642_620402# vssa1 0.41f
C1497 pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT vssa1 8.08f
C1498 a_343294_620745# vssa1 0.41f
C1499 pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN vssa1 12.9f
C1500 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT vssa1 13f
C1501 gpio_analog[3] vssa1 0.233p
C1502 a_339370_618592# vssa1 0.267f
C1503 io_out[11] vssa1 0.254p
C1504 a_339370_617808# vssa1 0.339f
C1505 a_336716_619863# vssa1 0.941f
C1506 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2 vssa1 9.9f
C1507 a_337674_622496# vssa1 0.267f
C1508 a_337674_621712# vssa1 0.311f
C1509 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1 vssa1 3.62f
C1510 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg vssa1 7.38f
C1511 io_out[15] vssa1 0.226p
C1512 w_336471_617254# vssa1 6.69f
C1513 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT vssa1 13.6f
C1514 vdda1 vssa1 0.742p
C1515 vccd1 vssa1 0.791p
C1516 io_out[12].t0 vssa1 0.173f
C1517 io_out[12].t1 vssa1 0.185f
C1518 io_out[12].n0 vssa1 1.18f
C1519 pmu_circuits_0.ldo_vb vssa1 38.3f
C1520 a_345642_614374.t4 vssa1 1.01f
C1521 a_345642_614374.t3 vssa1 0.946f
C1522 a_345642_614374.n0 vssa1 0.234f
C1523 a_345642_614374.t0 vssa1 0.451f
C1524 a_345642_614374.t2 vssa1 0.0858f
C1525 a_345642_614374.n1 vssa1 0.91f
C1526 a_345642_614374.n2 vssa1 0.154f
C1527 a_345642_614374.t1 vssa1 0.939f
C1528 a_345642_614374.t6 vssa1 1.01f
C1529 a_345642_614374.n3 vssa1 0.244f
C1530 a_345642_614374.n4 vssa1 0.172f
C1531 a_345642_614374.t5 vssa1 0.95f
C1532 a_345642_619372.t5 vssa1 0.939f
C1533 a_345642_619372.t3 vssa1 0.95f
C1534 a_345642_619372.t1 vssa1 1.01f
C1535 a_345642_619372.t2 vssa1 0.946f
C1536 a_345642_619372.n0 vssa1 0.234f
C1537 a_345642_619372.t0 vssa1 0.451f
C1538 a_345642_619372.t6 vssa1 0.0858f
C1539 a_345642_619372.n1 vssa1 0.91f
C1540 a_345642_619372.n2 vssa1 0.154f
C1541 a_345642_619372.n3 vssa1 0.172f
C1542 a_345642_619372.n4 vssa1 0.244f
C1543 a_345642_619372.t4 vssa1 1.01f
C1544 a_345642_621038.t3 vssa1 1.01f
C1545 a_345642_621038.t4 vssa1 0.95f
C1546 a_345642_621038.t1 vssa1 0.939f
C1547 a_345642_621038.t2 vssa1 1.01f
C1548 a_345642_621038.n0 vssa1 0.244f
C1549 a_345642_621038.n1 vssa1 0.172f
C1550 a_345642_621038.t6 vssa1 0.451f
C1551 a_345642_621038.t0 vssa1 0.0858f
C1552 a_345642_621038.n2 vssa1 0.91f
C1553 a_345642_621038.n3 vssa1 0.154f
C1554 a_345642_621038.n4 vssa1 0.234f
C1555 a_345642_621038.t5 vssa1 0.946f
C1556 a_336843_616061.t2 vssa1 0.845f
C1557 a_336843_616061.t0 vssa1 0.0037f
C1558 a_336843_616061.n0 vssa1 1.41f
C1559 a_336843_616061.t1 vssa1 0.0412f
C1560 a_341818_618261.t0 vssa1 0.451f
C1561 a_341818_618261.t5 vssa1 0.0858f
C1562 a_341818_618261.n0 vssa1 0.91f
C1563 a_341818_618261.t2 vssa1 1.01f
C1564 a_341818_618261.t3 vssa1 0.946f
C1565 a_341818_618261.n1 vssa1 0.234f
C1566 a_341818_618261.n2 vssa1 0.154f
C1567 a_341818_618261.t6 vssa1 0.939f
C1568 a_341818_618261.t1 vssa1 1.01f
C1569 a_341818_618261.n3 vssa1 0.244f
C1570 a_341818_618261.n4 vssa1 0.172f
C1571 a_341818_618261.t4 vssa1 0.95f
C1572 a_335719_622037.n0 vssa1 0.606f
C1573 a_335719_622037.t4 vssa1 0.00857f
C1574 a_335719_622037.t5 vssa1 0.0398f
C1575 a_335719_622037.n1 vssa1 0.702f
C1576 a_335719_622037.t1 vssa1 0.0133f
C1577 a_335719_622037.t8 vssa1 0.104f
C1578 a_335719_622037.n2 vssa1 0.125f
C1579 a_335719_622037.n3 vssa1 0.0654f
C1580 a_335719_622037.t0 vssa1 0.0633f
C1581 a_335719_622037.t7 vssa1 0.0633f
C1582 a_335719_622037.n4 vssa1 0.0962f
C1583 a_335719_622037.n5 vssa1 0.0792f
C1584 a_335719_622037.t6 vssa1 0.0633f
C1585 a_335719_622037.n6 vssa1 0.0962f
C1586 a_335719_622037.t9 vssa1 0.104f
C1587 a_335719_622037.n7 vssa1 0.125f
C1588 a_335719_622037.n8 vssa1 0.0654f
C1589 a_335719_622037.t2 vssa1 0.0633f
C1590 a_335719_622037.t3 vssa1 0.0168f
C1591 a_345642_617706.t4 vssa1 0.939f
C1592 a_345642_617706.t2 vssa1 0.95f
C1593 a_345642_617706.t1 vssa1 1.01f
C1594 a_345642_617706.t0 vssa1 0.946f
C1595 a_345642_617706.n0 vssa1 0.234f
C1596 a_345642_617706.t6 vssa1 0.451f
C1597 a_345642_617706.t5 vssa1 0.0858f
C1598 a_345642_617706.n1 vssa1 0.91f
C1599 a_345642_617706.n2 vssa1 0.154f
C1600 a_345642_617706.n3 vssa1 0.172f
C1601 a_345642_617706.n4 vssa1 0.244f
C1602 a_345642_617706.t3 vssa1 1.01f
C1603 a_341818_619927.t3 vssa1 1.02f
C1604 a_341818_619927.t4 vssa1 0.963f
C1605 a_341818_619927.t1 vssa1 0.952f
C1606 a_341818_619927.t2 vssa1 1.02f
C1607 a_341818_619927.n0 vssa1 0.247f
C1608 a_341818_619927.n1 vssa1 0.175f
C1609 a_341818_619927.t6 vssa1 0.458f
C1610 a_341818_619927.t0 vssa1 0.087f
C1611 a_341818_619927.n2 vssa1 0.923f
C1612 a_341818_619927.n3 vssa1 0.156f
C1613 a_341818_619927.n4 vssa1 0.238f
C1614 a_341818_619927.t5 vssa1 0.959f
C1615 io_out[11].t3 vssa1 0.00251f
C1616 io_out[11].t2 vssa1 0.00251f
C1617 io_out[11].n0 vssa1 0.0643f
C1618 pmu_circuits_0.iref_2nA_0.IREF vssa1 0.596f
C1619 io_out[11].t4 vssa1 0.0231f
C1620 pmu_circuits_0.vref01_0.VREF vssa1 4.65e-19
C1621 io_out[11].n1 vssa1 0.0233f
C1622 io_out[11].t1 vssa1 6.72e-19
C1623 io_out[11].t0 vssa1 0.00142f
C1624 io_out[11].n2 vssa1 0.0387f
C1625 io_out[11].n3 vssa1 0.067f
C1626 pmu_circuits_0.vref vssa1 2.3f
C1627 io_out[11].n4 vssa1 26.5f
C1628 pmu_circuits_0.iref vssa1 9.76f
C1629 a_352038_622652.n0 vssa1 0.342f
C1630 a_352038_622652.t0 vssa1 0.125f
C1631 a_352038_622652.t1 vssa1 0.0795f
C1632 a_352038_622652.n1 vssa1 0.291f
C1633 a_352038_622652.t2 vssa1 0.124f
C1634 a_352038_622652.n2 vssa1 0.157f
C1635 a_352038_622652.t6 vssa1 0.0336f
C1636 a_352038_622652.n3 vssa1 0.0907f
C1637 a_352038_622652.t4 vssa1 0.15f
C1638 a_352038_622652.n4 vssa1 0.278f
C1639 a_352038_622652.t5 vssa1 0.00593f
C1640 a_352038_622652.n5 vssa1 0.12f
C1641 a_352038_622652.n6 vssa1 0.239f
C1642 a_352038_622652.n7 vssa1 0.0463f
C1643 a_352038_622652.t3 vssa1 0.0185f
C1644 io_out[15].t4 vssa1 0.00907f
C1645 io_out[15].n0 vssa1 0.00588f
C1646 io_out[15].t1 vssa1 0.0578f
C1647 io_out[15].n1 vssa1 0.116f
C1648 io_out[15].n2 vssa1 0.0109f
C1649 io_out[15].n3 vssa1 0.0218f
C1650 io_out[15].n4 vssa1 0.00393f
C1651 io_out[15].n5 vssa1 0.202f
C1652 io_out[15].n6 vssa1 0.0253f
C1653 io_out[15].n7 vssa1 0.0253f
C1654 io_out[15].n8 vssa1 0.0214f
C1655 io_out[15].n9 vssa1 0.183f
C1656 io_out[15].n10 vssa1 0.261f
C1657 io_out[15].n11 vssa1 0.0122f
C1658 io_out[15].n13 vssa1 0.00392f
C1659 io_out[15].n14 vssa1 0.153f
C1660 io_out[15].t0 vssa1 0.0182f
C1661 io_out[15].n15 vssa1 0.139f
C1662 io_out[15].n16 vssa1 0.28f
C1663 io_out[15].n17 vssa1 0.0127f
C1664 io_out[15].n18 vssa1 0.0114f
C1665 io_out[15].t2 vssa1 0.00935f
C1666 io_out[15].n19 vssa1 0.0397f
C1667 io_out[15].n20 vssa1 0.0201f
C1668 io_out[15].n21 vssa1 0.00491f
C1669 io_out[15].n22 vssa1 0.00785f
C1670 io_out[15].n23 vssa1 0.0474f
C1671 io_out[15].t3 vssa1 2.3f
C1672 io_out[15].n24 vssa1 0.171f
C1673 pmu_circuits_0.ldo_out vssa1 0.0465f
C1674 io_out[15].n25 vssa1 24f
C1675 io_out[16].t0 vssa1 0.0919f
C1676 io_out[16].t1 vssa1 0.114f
C1677 io_out[16].n0 vssa1 8.31e-20
C1678 pmu_circuits_0.ldo_vs vssa1 0.00337f
C1679 io_out[16].n1 vssa1 15f
C1680 a_345642_616040.t3 vssa1 0.946f
C1681 a_345642_616040.t2 vssa1 0.95f
C1682 a_345642_616040.t1 vssa1 0.939f
C1683 a_345642_616040.t4 vssa1 1.01f
C1684 a_345642_616040.n0 vssa1 0.244f
C1685 a_345642_616040.n1 vssa1 0.172f
C1686 a_345642_616040.t6 vssa1 0.451f
C1687 a_345642_616040.t0 vssa1 0.0858f
C1688 a_345642_616040.n2 vssa1 0.91f
C1689 a_345642_616040.n3 vssa1 0.154f
C1690 a_345642_616040.n4 vssa1 0.234f
C1691 a_345642_616040.t5 vssa1 1.01f
C1692 a_341818_613263.t1 vssa1 0.939f
C1693 a_341818_613263.t4 vssa1 0.95f
C1694 a_341818_613263.t6 vssa1 0.451f
C1695 a_341818_613263.t0 vssa1 0.0858f
C1696 a_341818_613263.n0 vssa1 0.91f
C1697 a_341818_613263.t3 vssa1 1.01f
C1698 a_341818_613263.t2 vssa1 0.946f
C1699 a_341818_613263.n1 vssa1 0.234f
C1700 a_341818_613263.n2 vssa1 0.154f
C1701 a_341818_613263.n3 vssa1 0.172f
C1702 a_341818_613263.n4 vssa1 0.244f
C1703 a_341818_613263.t5 vssa1 1.01f
C1704 pmu_circuits_0.ring_100mV_0.mdls_inv_1.IN vssa1 0.484f
C1705 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n0 vssa1 0.299f
C1706 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n1 vssa1 0.312f
C1707 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t2 vssa1 0.652f
C1708 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t4 vssa1 0.652f
C1709 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t0 vssa1 0.696f
C1710 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n2 vssa1 0.194f
C1711 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n3 vssa1 0.186f
C1712 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t3 vssa1 0.0589f
C1713 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n4 vssa1 0.494f
C1714 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t11 vssa1 0.181f
C1715 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t7 vssa1 0.182f
C1716 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n5 vssa1 0.529f
C1717 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t14 vssa1 0.233f
C1718 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n6 vssa1 0.0909f
C1719 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n7 vssa1 0.448f
C1720 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n8 vssa1 0.58f
C1721 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t9 vssa1 0.36f
C1722 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t10 vssa1 0.357f
C1723 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n9 vssa1 0.582f
C1724 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t5 vssa1 0.358f
C1725 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n10 vssa1 0.582f
C1726 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t8 vssa1 0.357f
C1727 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t12 vssa1 0.448f
C1728 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n11 vssa1 0.351f
C1729 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n12 vssa1 0.117f
C1730 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n13 vssa1 0.35f
C1731 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t6 vssa1 0.447f
C1732 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n14 vssa1 0.335f
C1733 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t15 vssa1 0.482f
C1734 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n15 vssa1 0.801f
C1735 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n16 vssa1 0.847f
C1736 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t13 vssa1 0.166f
C1737 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.t1 vssa1 0.0107f
C1738 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n17 vssa1 0.123f
C1739 pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT.n18 vssa1 0.315f
C1740 a_350722_615130.t7 vssa1 0.0645f
C1741 a_350722_615130.t5 vssa1 0.0644f
C1742 a_350722_615130.t4 vssa1 0.0716f
C1743 a_350722_615130.t0 vssa1 0.144f
C1744 a_350722_615130.t3 vssa1 0.0219f
C1745 a_350722_615130.n0 vssa1 0.546f
C1746 a_350722_615130.n1 vssa1 0.418f
C1747 a_350722_615130.n2 vssa1 0.243f
C1748 a_350722_615130.n3 vssa1 0.243f
C1749 a_350722_615130.t1 vssa1 0.0908f
C1750 a_350722_615130.t2 vssa1 0.0757f
C1751 a_350722_615130.n4 vssa1 0.875f
C1752 a_350722_615130.n5 vssa1 0.471f
C1753 a_350722_615130.t6 vssa1 0.0714f
C1754 gpio_analog[7].n0 vssa1 0.0131f
C1755 gpio_analog[7].t0 vssa1 0.0149f
C1756 gpio_analog[7].n1 vssa1 0.0131f
C1757 gpio_analog[7].t4 vssa1 0.0149f
C1758 gpio_analog[7].n2 vssa1 0.0207f
C1759 gpio_analog[7].t5 vssa1 0.0149f
C1760 gpio_analog[7].t9 vssa1 0.0196f
C1761 gpio_analog[7].n3 vssa1 0.0294f
C1762 gpio_analog[7].n4 vssa1 0.0157f
C1763 gpio_analog[7].n5 vssa1 0.0138f
C1764 gpio_analog[7].t7 vssa1 0.0196f
C1765 gpio_analog[7].n6 vssa1 0.0207f
C1766 gpio_analog[7].t8 vssa1 0.0149f
C1767 gpio_analog[7].n7 vssa1 0.0294f
C1768 gpio_analog[7].n8 vssa1 0.0131f
C1769 gpio_analog[7].t6 vssa1 0.0149f
C1770 gpio_analog[7].n9 vssa1 0.0157f
C1771 gpio_analog[7].n10 vssa1 0.0131f
C1772 gpio_analog[7].t2 vssa1 0.0149f
C1773 gpio_analog[7].n11 vssa1 0.0137f
C1774 gpio_analog[7].t1 vssa1 0.00296f
C1775 gpio_analog[7].t3 vssa1 0.00296f
C1776 gpio_analog[7].n12 vssa1 0.0675f
C1777 gpio_analog[7].n13 vssa1 0.0465f
C1778 pmu_circuits_0.ldo_iref vssa1 6.5f
C1779 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t12 vssa1 0.153f
C1780 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t15 vssa1 0.152f
C1781 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n0 vssa1 0.445f
C1782 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t14 vssa1 0.196f
C1783 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n1 vssa1 0.0764f
C1784 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n2 vssa1 0.377f
C1785 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n3 vssa1 0.251f
C1786 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n4 vssa1 0.488f
C1787 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t10 vssa1 0.302f
C1788 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t7 vssa1 0.3f
C1789 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n5 vssa1 0.489f
C1790 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t13 vssa1 0.301f
C1791 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n6 vssa1 0.489f
C1792 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t6 vssa1 0.3f
C1793 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n7 vssa1 0.227f
C1794 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n8 vssa1 0.0354f
C1795 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t11 vssa1 0.376f
C1796 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n9 vssa1 0.296f
C1797 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n10 vssa1 0.0983f
C1798 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n11 vssa1 0.294f
C1799 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t8 vssa1 0.376f
C1800 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n12 vssa1 0.307f
C1801 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n13 vssa1 0.282f
C1802 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t5 vssa1 0.406f
C1803 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n14 vssa1 0.64f
C1804 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n15 vssa1 0.605f
C1805 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t9 vssa1 0.14f
C1806 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t4 vssa1 0.009f
C1807 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n16 vssa1 0.103f
C1808 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n17 vssa1 0.265f
C1809 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n18 vssa1 0.376f
C1810 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t2 vssa1 0.548f
C1811 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t0 vssa1 0.548f
C1812 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t1 vssa1 0.585f
C1813 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n19 vssa1 0.163f
C1814 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n20 vssa1 0.157f
C1815 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.t3 vssa1 0.0495f
C1816 pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN.n21 vssa1 0.412f
C1817 pmu_circuits_0.ring_100mV_0.mdls_inv_6.OUT vssa1 0.0825f
C1818 a_341818_616595.t6 vssa1 0.458f
C1819 a_341818_616595.t2 vssa1 0.963f
C1820 a_341818_616595.t0 vssa1 0.952f
C1821 a_341818_616595.t3 vssa1 1.02f
C1822 a_341818_616595.n0 vssa1 0.247f
C1823 a_341818_616595.n1 vssa1 0.175f
C1824 a_341818_616595.t5 vssa1 1.02f
C1825 a_341818_616595.t4 vssa1 0.959f
C1826 a_341818_616595.n2 vssa1 0.238f
C1827 a_341818_616595.n3 vssa1 0.156f
C1828 a_341818_616595.n4 vssa1 0.923f
C1829 a_341818_616595.t1 vssa1 0.087f
C1830 a_341818_614929.t0 vssa1 0.939f
C1831 a_341818_614929.t3 vssa1 0.95f
C1832 a_341818_614929.t6 vssa1 0.451f
C1833 a_341818_614929.t1 vssa1 0.0858f
C1834 a_341818_614929.n0 vssa1 0.91f
C1835 a_341818_614929.t2 vssa1 1.01f
C1836 a_341818_614929.t4 vssa1 0.946f
C1837 a_341818_614929.n1 vssa1 0.234f
C1838 a_341818_614929.n2 vssa1 0.154f
C1839 a_341818_614929.n3 vssa1 0.172f
C1840 a_341818_614929.n4 vssa1 0.244f
C1841 a_341818_614929.t5 vssa1 1.01f
C1842 pmu_circuits_0.ring_100mV_0.mdls_inv_8.IN vssa1 0.407f
C1843 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n0 vssa1 0.251f
C1844 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n1 vssa1 0.263f
C1845 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t15 vssa1 0.153f
C1846 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t6 vssa1 0.152f
C1847 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n2 vssa1 0.445f
C1848 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t12 vssa1 0.196f
C1849 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n3 vssa1 0.0764f
C1850 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n4 vssa1 0.377f
C1851 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n5 vssa1 0.488f
C1852 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t14 vssa1 0.302f
C1853 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t9 vssa1 0.3f
C1854 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n6 vssa1 0.489f
C1855 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t7 vssa1 0.301f
C1856 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n7 vssa1 0.489f
C1857 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t11 vssa1 0.3f
C1858 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t5 vssa1 0.376f
C1859 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n8 vssa1 0.295f
C1860 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n9 vssa1 0.0983f
C1861 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n10 vssa1 0.294f
C1862 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t10 vssa1 0.376f
C1863 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n11 vssa1 0.282f
C1864 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t8 vssa1 0.406f
C1865 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n12 vssa1 0.641f
C1866 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n13 vssa1 0.606f
C1867 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t13 vssa1 0.14f
C1868 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t0 vssa1 0.009f
C1869 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n14 vssa1 0.103f
C1870 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n15 vssa1 0.265f
C1871 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n16 vssa1 0.376f
C1872 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t2 vssa1 0.548f
C1873 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t4 vssa1 0.585f
C1874 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n17 vssa1 0.163f
C1875 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t1 vssa1 0.548f
C1876 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n18 vssa1 0.157f
C1877 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.t3 vssa1 0.0495f
C1878 pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT.n19 vssa1 0.412f
C1879 pmu_circuits_0.ring_out vssa1 0.00203f
C1880 gpio_analog[3].t19 vssa1 0.00255f
C1881 gpio_analog[3].t16 vssa1 0.00171f
C1882 gpio_analog[3].n0 vssa1 0.0485f
C1883 gpio_analog[3].t17 vssa1 0.00171f
C1884 gpio_analog[3].n1 vssa1 0.0253f
C1885 gpio_analog[3].t18 vssa1 0.00204f
C1886 gpio_analog[3].n2 vssa1 0.0282f
C1887 gpio_analog[3].t12 vssa1 0.03f
C1888 gpio_analog[3].n3 vssa1 0.0229f
C1889 gpio_analog[3].t10 vssa1 0.0296f
C1890 gpio_analog[3].t1 vssa1 0.0296f
C1891 gpio_analog[3].t0 vssa1 0.0457f
C1892 gpio_analog[3].t9 vssa1 0.0303f
C1893 gpio_analog[3].n4 vssa1 0.12f
C1894 gpio_analog[3].t11 vssa1 0.0303f
C1895 gpio_analog[3].n5 vssa1 0.0692f
C1896 gpio_analog[3].t13 vssa1 0.0303f
C1897 gpio_analog[3].n6 vssa1 0.0692f
C1898 gpio_analog[3].t7 vssa1 0.0303f
C1899 gpio_analog[3].n7 vssa1 0.0692f
C1900 gpio_analog[3].t8 vssa1 0.0303f
C1901 gpio_analog[3].n8 vssa1 0.0692f
C1902 gpio_analog[3].t4 vssa1 0.0303f
C1903 gpio_analog[3].n9 vssa1 0.0692f
C1904 gpio_analog[3].t5 vssa1 0.0303f
C1905 gpio_analog[3].n10 vssa1 0.0692f
C1906 gpio_analog[3].t6 vssa1 0.0303f
C1907 gpio_analog[3].n11 vssa1 0.0692f
C1908 gpio_analog[3].t2 vssa1 0.0303f
C1909 gpio_analog[3].n12 vssa1 0.0692f
C1910 gpio_analog[3].t3 vssa1 0.0303f
C1911 gpio_analog[3].n13 vssa1 0.0692f
C1912 gpio_analog[3].t14 vssa1 0.0303f
C1913 gpio_analog[3].n14 vssa1 0.0692f
C1914 gpio_analog[3].t15 vssa1 0.0303f
C1915 gpio_analog[3].n15 vssa1 0.0699f
C1916 gpio_analog[3].n16 vssa1 0.124f
C1917 gpio_analog[3].n17 vssa1 0.0951f
C1918 gpio_analog[3].n18 vssa1 0.279f
C1919 gpio_analog[3].n19 vssa1 19.2f
C1920 a_341600_622217.t3 vssa1 0.205f
C1921 a_341600_622217.t0 vssa1 0.139f
C1922 a_341600_622217.n0 vssa1 0.527f
C1923 a_341600_622217.t1 vssa1 0.139f
C1924 a_341600_622217.n1 vssa1 0.303f
C1925 a_341600_622217.t2 vssa1 0.139f
C1926 a_341600_622217.n2 vssa1 0.303f
C1927 a_341600_622217.t6 vssa1 0.139f
C1928 a_341600_622217.n3 vssa1 0.303f
C1929 a_341600_622217.t29 vssa1 0.194f
C1930 a_341600_622217.n4 vssa1 0.251f
C1931 a_341600_622217.t19 vssa1 0.194f
C1932 a_341600_622217.n5 vssa1 0.263f
C1933 a_341600_622217.t16 vssa1 0.194f
C1934 a_341600_622217.n6 vssa1 0.149f
C1935 a_341600_622217.t13 vssa1 0.194f
C1936 a_341600_622217.n7 vssa1 0.149f
C1937 a_341600_622217.t21 vssa1 0.194f
C1938 a_341600_622217.n8 vssa1 0.149f
C1939 a_341600_622217.t20 vssa1 0.194f
C1940 a_341600_622217.n9 vssa1 0.149f
C1941 a_341600_622217.n10 vssa1 0.267f
C1942 a_341600_622217.n11 vssa1 0.149f
C1943 a_341600_622217.n12 vssa1 0.149f
C1944 a_341600_622217.n13 vssa1 0.149f
C1945 a_341600_622217.n14 vssa1 0.149f
C1946 a_341600_622217.n15 vssa1 0.149f
C1947 a_341600_622217.t24 vssa1 0.194f
C1948 a_341600_622217.n16 vssa1 0.149f
C1949 a_341600_622217.t23 vssa1 0.194f
C1950 a_341600_622217.n17 vssa1 0.149f
C1951 a_341600_622217.n18 vssa1 0.149f
C1952 a_341600_622217.n19 vssa1 0.149f
C1953 a_341600_622217.t22 vssa1 0.194f
C1954 a_341600_622217.n20 vssa1 0.149f
C1955 a_341600_622217.t26 vssa1 0.194f
C1956 a_341600_622217.n21 vssa1 0.149f
C1957 a_341600_622217.n22 vssa1 0.149f
C1958 a_341600_622217.n23 vssa1 0.149f
C1959 a_341600_622217.t25 vssa1 0.194f
C1960 a_341600_622217.n24 vssa1 0.139f
C1961 a_341600_622217.t14 vssa1 0.322f
C1962 a_341600_622217.t17 vssa1 0.194f
C1963 a_341600_622217.n25 vssa1 0.226f
C1964 a_341600_622217.t27 vssa1 0.194f
C1965 a_341600_622217.n26 vssa1 0.149f
C1966 a_341600_622217.t10 vssa1 0.194f
C1967 a_341600_622217.n27 vssa1 0.149f
C1968 a_341600_622217.n28 vssa1 0.226f
C1969 a_341600_622217.n29 vssa1 0.149f
C1970 a_341600_622217.n30 vssa1 0.149f
C1971 a_341600_622217.n31 vssa1 0.149f
C1972 a_341600_622217.t12 vssa1 0.194f
C1973 a_341600_622217.n32 vssa1 0.14f
C1974 a_341600_622217.n33 vssa1 0.104f
C1975 a_341600_622217.t9 vssa1 0.00583f
C1976 a_341600_622217.t15 vssa1 0.125f
C1977 a_341600_622217.n34 vssa1 0.0749f
C1978 a_341600_622217.t18 vssa1 0.0527f
C1979 a_341600_622217.n35 vssa1 0.0889f
C1980 a_341600_622217.t28 vssa1 0.0527f
C1981 a_341600_622217.n36 vssa1 0.0707f
C1982 a_341600_622217.n37 vssa1 0.0889f
C1983 a_341600_622217.n38 vssa1 0.0707f
C1984 a_341600_622217.n39 vssa1 0.0561f
C1985 a_341600_622217.n40 vssa1 0.0295f
C1986 a_341600_622217.t11 vssa1 0.0885f
C1987 a_341600_622217.n41 vssa1 0.0928f
C1988 a_341600_622217.n42 vssa1 0.139f
C1989 a_341600_622217.t8 vssa1 0.011f
C1990 a_341600_622217.n43 vssa1 0.568f
C1991 a_341600_622217.t5 vssa1 0.139f
C1992 a_341600_622217.n44 vssa1 0.327f
C1993 a_341600_622217.t4 vssa1 0.139f
C1994 a_341600_622217.n45 vssa1 0.303f
C1995 a_341600_622217.n46 vssa1 0.303f
C1996 a_341600_622217.t7 vssa1 0.139f
C1997 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n0 vssa1 1.59f
C1998 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t15 vssa1 0.13f
C1999 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t8 vssa1 0.129f
C2000 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n1 vssa1 0.378f
C2001 pmu_circuits_0.ring_100mV_0.ring_100mV_buffer_0.IN vssa1 0.443f
C2002 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t13 vssa1 0.164f
C2003 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t16 vssa1 0.176f
C2004 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n2 vssa1 0.0691f
C2005 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n3 vssa1 0.387f
C2006 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n4 vssa1 0.235f
C2007 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n5 vssa1 0.235f
C2008 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n6 vssa1 0.235f
C2009 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n7 vssa1 0.235f
C2010 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n8 vssa1 0.235f
C2011 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n9 vssa1 0.306f
C2012 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t7 vssa1 0.255f
C2013 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t5 vssa1 0.255f
C2014 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t12 vssa1 0.255f
C2015 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t17 vssa1 0.255f
C2016 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t10 vssa1 0.374f
C2017 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n10 vssa1 0.393f
C2018 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t14 vssa1 0.255f
C2019 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n11 vssa1 0.238f
C2020 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n12 vssa1 0.238f
C2021 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t6 vssa1 0.255f
C2022 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n13 vssa1 0.238f
C2023 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n14 vssa1 0.238f
C2024 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t9 vssa1 0.255f
C2025 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n15 vssa1 0.238f
C2026 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n16 vssa1 0.224f
C2027 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n17 vssa1 0.151f
C2028 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n18 vssa1 0.529f
C2029 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t11 vssa1 0.118f
C2030 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t4 vssa1 0.00764f
C2031 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n19 vssa1 0.0878f
C2032 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n20 vssa1 0.225f
C2033 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n21 vssa1 0.319f
C2034 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t3 vssa1 0.465f
C2035 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t2 vssa1 0.465f
C2036 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t0 vssa1 0.496f
C2037 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n22 vssa1 0.138f
C2038 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n23 vssa1 0.133f
C2039 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.t1 vssa1 0.042f
C2040 pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT.n24 vssa1 0.35f
C2041 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n0 vssa1 0.249f
C2042 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n1 vssa1 0.261f
C2043 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t8 vssa1 0.151f
C2044 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t11 vssa1 0.151f
C2045 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n2 vssa1 0.441f
C2046 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t10 vssa1 0.194f
C2047 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n3 vssa1 0.0758f
C2048 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n4 vssa1 0.374f
C2049 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n5 vssa1 0.484f
C2050 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t6 vssa1 0.3f
C2051 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t7 vssa1 0.298f
C2052 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n6 vssa1 0.485f
C2053 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t12 vssa1 0.299f
C2054 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n7 vssa1 0.485f
C2055 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t14 vssa1 0.298f
C2056 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t9 vssa1 0.373f
C2057 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n8 vssa1 0.293f
C2058 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n9 vssa1 0.0975f
C2059 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n10 vssa1 0.292f
C2060 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t13 vssa1 0.373f
C2061 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n11 vssa1 0.279f
C2062 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t5 vssa1 0.402f
C2063 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n12 vssa1 0.636f
C2064 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n13 vssa1 0.594f
C2065 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t15 vssa1 0.138f
C2066 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t2 vssa1 0.00893f
C2067 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n14 vssa1 0.103f
C2068 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n15 vssa1 0.263f
C2069 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n16 vssa1 0.373f
C2070 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t1 vssa1 0.544f
C2071 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t4 vssa1 0.58f
C2072 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t0 vssa1 0.544f
C2073 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n17 vssa1 0.162f
C2074 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n18 vssa1 0.155f
C2075 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.t3 vssa1 0.0491f
C2076 pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN.n19 vssa1 0.409f
C2077 pmu_circuits_0.ring_100mV_0.mdls_inv_8.OUT vssa1 0.0818f
C2078 pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Ip1 vssa1 0.953f
C2079 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t0 vssa1 0.0634f
C2080 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t2 vssa1 0.0268f
C2081 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t3 vssa1 0.0271f
C2082 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t6 vssa1 0.557f
C2083 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t5 vssa1 0.453f
C2084 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n0 vssa1 1.59f
C2085 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t4 vssa1 0.453f
C2086 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n1 vssa1 0.852f
C2087 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t7 vssa1 0.453f
C2088 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n2 vssa1 0.977f
C2089 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n3 vssa1 0.838f
C2090 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.n4 vssa1 0.721f
C2091 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1.t1 vssa1 0.0364f
C2092 a_350378_615130.n0 vssa1 0.797f
C2093 a_350378_615130.t4 vssa1 0.069f
C2094 a_350378_615130.t3 vssa1 0.00829f
C2095 a_350378_615130.t2 vssa1 0.00528f
C2096 a_350378_615130.t5 vssa1 6.57f
C2097 a_350378_615130.n1 vssa1 1.14f
C2098 a_350378_615130.t1 vssa1 0.0995f
C2099 a_350378_615130.n2 vssa1 0.889f
C2100 a_350378_615130.t0 vssa1 0.0229f
C2101 a_350942_613328.n0 vssa1 1.03f
C2102 a_350942_613328.t5 vssa1 0.351f
C2103 a_350942_613328.t7 vssa1 0.719f
C2104 a_350942_613328.t2 vssa1 0.429f
C2105 a_350942_613328.n1 vssa1 0.229f
C2106 a_350942_613328.t3 vssa1 0.00554f
C2107 a_350942_613328.t6 vssa1 0.719f
C2108 a_350942_613328.t0 vssa1 0.429f
C2109 a_350942_613328.n2 vssa1 0.229f
C2110 a_350942_613328.t1 vssa1 0.00554f
C2111 a_350942_613328.n3 vssa1 1.09f
C2112 a_350942_613328.t4 vssa1 0.162f
C2113 a_339370_613888.n0 vssa1 0.9f
C2114 a_339370_613888.n1 vssa1 0.9f
C2115 a_339370_613888.t16 vssa1 0.028f
C2116 a_339370_613888.t7 vssa1 0.0279f
C2117 a_339370_613888.n2 vssa1 0.372f
C2118 a_339370_613888.t14 vssa1 0.028f
C2119 a_339370_613888.t5 vssa1 0.0279f
C2120 a_339370_613888.n3 vssa1 0.45f
C2121 a_339370_613888.t13 vssa1 0.028f
C2122 a_339370_613888.t4 vssa1 0.0279f
C2123 a_339370_613888.n4 vssa1 0.45f
C2124 a_339370_613888.t11 vssa1 0.028f
C2125 a_339370_613888.t2 vssa1 0.0279f
C2126 a_339370_613888.n5 vssa1 0.448f
C2127 a_339370_613888.t19 vssa1 0.028f
C2128 a_339370_613888.t0 vssa1 0.0279f
C2129 a_339370_613888.t15 vssa1 0.028f
C2130 a_339370_613888.t6 vssa1 0.0279f
C2131 a_339370_613888.n6 vssa1 0.372f
C2132 a_339370_613888.t17 vssa1 0.028f
C2133 a_339370_613888.t8 vssa1 0.0279f
C2134 a_339370_613888.n7 vssa1 0.45f
C2135 a_339370_613888.t10 vssa1 0.028f
C2136 a_339370_613888.t1 vssa1 0.0279f
C2137 a_339370_613888.n8 vssa1 0.45f
C2138 a_339370_613888.t12 vssa1 0.028f
C2139 a_339370_613888.t3 vssa1 0.0279f
C2140 a_339370_613888.n9 vssa1 0.448f
C2141 a_339370_613888.t18 vssa1 0.028f
C2142 a_339370_613888.t9 vssa1 0.0279f
C2143 pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Ip2 vssa1 1.97f
C2144 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n0 vssa1 0.694f
C2145 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n1 vssa1 1.36f
C2146 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t3 vssa1 0.0454f
C2147 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t11 vssa1 0.0194f
C2148 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n2 vssa1 0.562f
C2149 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t10 vssa1 0.0194f
C2150 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t7 vssa1 0.0194f
C2151 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t8 vssa1 0.0454f
C2152 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n3 vssa1 0.561f
C2153 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t5 vssa1 0.0454f
C2154 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t9 vssa1 0.0194f
C2155 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n4 vssa1 0.562f
C2156 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t6 vssa1 0.0194f
C2157 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t4 vssa1 0.0194f
C2158 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t2 vssa1 0.0454f
C2159 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n5 vssa1 0.561f
C2160 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t15 vssa1 0.971f
C2161 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t18 vssa1 1.03f
C2162 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t19 vssa1 1.03f
C2163 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t23 vssa1 1.03f
C2164 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t13 vssa1 1.03f
C2165 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t22 vssa1 1.03f
C2166 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t16 vssa1 1.03f
C2167 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t24 vssa1 1.03f
C2168 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t21 vssa1 1.03f
C2169 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t12 vssa1 1.03f
C2170 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t20 vssa1 1.03f
C2171 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t25 vssa1 1.03f
C2172 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t14 vssa1 0.683f
C2173 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t17 vssa1 0.625f
C2174 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n6 vssa1 1.14f
C2175 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t0 vssa1 0.0407f
C2176 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.n7 vssa1 0.956f
C2177 pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2.t1 vssa1 0.0281f
C2178 a_335807_622237.n0 vssa1 0.705f
C2179 a_335807_622237.n1 vssa1 3.28f
C2180 a_335807_622237.t1 vssa1 0.0167f
C2181 a_335807_622237.t7 vssa1 0.888f
C2182 a_335807_622237.t15 vssa1 0.902f
C2183 a_335807_622237.t21 vssa1 0.828f
C2184 a_335807_622237.t22 vssa1 0.475f
C2185 a_335807_622237.n2 vssa1 0.799f
C2186 a_335807_622237.t9 vssa1 1.62f
C2187 a_335807_622237.t12 vssa1 0.887f
C2188 a_335807_622237.t13 vssa1 0.887f
C2189 a_335807_622237.t18 vssa1 0.887f
C2190 a_335807_622237.t6 vssa1 0.887f
C2191 a_335807_622237.t17 vssa1 0.887f
C2192 a_335807_622237.t10 vssa1 0.887f
C2193 a_335807_622237.t19 vssa1 0.887f
C2194 a_335807_622237.t16 vssa1 0.887f
C2195 a_335807_622237.t23 vssa1 0.887f
C2196 a_335807_622237.t14 vssa1 0.887f
C2197 a_335807_622237.t20 vssa1 0.887f
C2198 a_335807_622237.t8 vssa1 0.887f
C2199 a_335807_622237.t11 vssa1 0.627f
C2200 a_335807_622237.t4 vssa1 0.126f
C2201 a_335807_622237.t5 vssa1 0.218f
C2202 a_335807_622237.n3 vssa1 2.68f
C2203 a_335807_622237.n4 vssa1 0.151f
C2204 a_335807_622237.t2 vssa1 0.298f
C2205 a_335807_622237.t0 vssa1 0.294f
C2206 a_335807_622237.n5 vssa1 0.432f
C2207 a_335807_622237.t3 vssa1 0.0167f
C2208 VCCD1 vssa1 2.53f
C2209 vccd1.n0 vssa1 46.4f
C2210 vccd1.t58 vssa1 0.00191f
C2211 vccd1.t59 vssa1 0.00235f
C2212 pmu_circuits_0.vref01_0.DD vssa1 0.00469f
C2213 vccd1.n1 vssa1 0.00466f
C2214 vccd1.t54 vssa1 0.00367f
C2215 vccd1.n2 vssa1 0.00394f
C2216 vccd1.n3 vssa1 1.17e-19
C2217 vccd1.n4 vssa1 6.69e-19
C2218 vccd1.n5 vssa1 4.68e-19
C2219 vccd1.n6 vssa1 7.11e-19
C2220 vccd1.n7 vssa1 0.00103f
C2221 vccd1.n8 vssa1 0.0193f
C2222 vccd1.n9 vssa1 0.0103f
C2223 vccd1.t31 vssa1 0.00784f
C2224 vccd1.n10 vssa1 0.00493f
C2225 vccd1.n11 vssa1 7.28e-19
C2226 vccd1.n12 vssa1 8.2e-19
C2227 vccd1.t49 vssa1 4.42e-19
C2228 vccd1.n14 vssa1 0.00629f
C2229 vccd1.n15 vssa1 8.53e-19
C2230 vccd1.n16 vssa1 8.53e-19
C2231 vccd1.t48 vssa1 0.00937f
C2232 vccd1.n18 vssa1 0.00629f
C2233 vccd1.n19 vssa1 8.53e-19
C2234 vccd1.n20 vssa1 0.0035f
C2235 vccd1.n21 vssa1 0.0026f
C2236 vccd1.t13 vssa1 3.6e-19
C2237 vccd1.n22 vssa1 0.00155f
C2238 vccd1.n23 vssa1 0.0102f
C2239 vccd1.t32 vssa1 0.0156f
C2240 vccd1.t67 vssa1 0.019f
C2241 vccd1.t46 vssa1 0.014f
C2242 vccd1.n24 vssa1 0.00952f
C2243 vccd1.n25 vssa1 0.00214f
C2244 vccd1.t33 vssa1 2.28e-19
C2245 vccd1.n26 vssa1 0.00229f
C2246 vccd1.t68 vssa1 7.6e-20
C2247 vccd1.n27 vssa1 0.00303f
C2248 vccd1.t47 vssa1 7.6e-20
C2249 vccd1.n28 vssa1 0.00257f
C2250 vccd1.n29 vssa1 0.00127f
C2251 vccd1.t45 vssa1 7.6e-20
C2252 vccd1.n30 vssa1 0.00264f
C2253 vccd1.t66 vssa1 7.6e-20
C2254 vccd1.n31 vssa1 0.00303f
C2255 vccd1.t12 vssa1 3.64e-19
C2256 vccd1.n32 vssa1 0.00232f
C2257 vccd1.t10 vssa1 0.00784f
C2258 vccd1.n33 vssa1 0.00662f
C2259 vccd1.t44 vssa1 0.0145f
C2260 vccd1.t65 vssa1 0.019f
C2261 vccd1.t11 vssa1 0.015f
C2262 vccd1.n34 vssa1 0.00969f
C2263 vccd1.n35 vssa1 0.00214f
C2264 vccd1.n36 vssa1 0.00121f
C2265 vccd1.t34 vssa1 3.6e-19
C2266 vccd1.n37 vssa1 0.00141f
C2267 vccd1.n38 vssa1 0.0085f
C2268 vccd1.n39 vssa1 0.00384f
C2269 vccd1.n40 vssa1 0.0143f
C2270 pmu_circuits_0.ldo_0.DD vssa1 0.0344f
C2271 vccd1.n41 vssa1 0.118f
C2272 vccd1.t56 vssa1 7.31e-19
C2273 vccd1.n42 vssa1 0.00465f
C2274 vccd1.n43 vssa1 0.0031f
C2275 vccd1.n44 vssa1 6.62e-19
C2276 vccd1.n45 vssa1 0.00894f
C2277 vccd1.n46 vssa1 0.0013f
C2278 vccd1.n47 vssa1 6.84e-19
C2279 vccd1.t1 vssa1 2.02e-19
C2280 vccd1.n48 vssa1 0.00216f
C2281 vccd1.n49 vssa1 0.00168f
C2282 vccd1.n50 vssa1 0.0148f
C2283 vccd1.n51 vssa1 0.0123f
C2284 vccd1.t15 vssa1 0.0117f
C2285 vccd1.t0 vssa1 0.00998f
C2286 vccd1.t43 vssa1 0.021f
C2287 vccd1.t14 vssa1 0.00395f
C2288 vccd1.t16 vssa1 4.27e-20
C2289 vccd1.n52 vssa1 0.00731f
C2290 vccd1.n53 vssa1 2.54e-19
C2291 vccd1.n54 vssa1 9.18e-19
C2292 vccd1.n55 vssa1 0.00146f
C2293 vccd1.n56 vssa1 0.00167f
C2294 vccd1.n57 vssa1 0.0218f
C2295 vccd1.n58 vssa1 0.00167f
C2296 vccd1.n59 vssa1 0.00109f
C2297 vccd1.n60 vssa1 0.0107f
C2298 vccd1.n61 vssa1 0.00665f
C2299 vccd1.n62 vssa1 0.00665f
C2300 vccd1.n63 vssa1 0.122f
C2301 vccd1.t21 vssa1 0.048f
C2302 vccd1.n64 vssa1 0.0028f
C2303 vccd1.n65 vssa1 0.0028f
C2304 vccd1.t75 vssa1 9.71e-19
C2305 vccd1.t64 vssa1 9.71e-19
C2306 vccd1.n66 vssa1 0.00144f
C2307 vccd1.n67 vssa1 0.00138f
C2308 vccd1.t22 vssa1 4.27e-20
C2309 vccd1.n68 vssa1 5.47e-19
C2310 vccd1.t8 vssa1 4.27e-20
C2311 vccd1.n69 vssa1 5.47e-19
C2312 vccd1.t19 vssa1 4.27e-20
C2313 vccd1.n70 vssa1 5.47e-19
C2314 vccd1.t37 vssa1 4.27e-20
C2315 vccd1.n71 vssa1 5.47e-19
C2316 vccd1.t51 vssa1 9.31e-19
C2317 vccd1.t60 vssa1 9.31e-19
C2318 vccd1.t61 vssa1 9.31e-19
C2319 vccd1.t74 vssa1 9.31e-19
C2320 vccd1.t70 vssa1 9.31e-19
C2321 vccd1.t73 vssa1 9.31e-19
C2322 vccd1.t52 vssa1 9.31e-19
C2323 vccd1.t41 vssa1 9.31e-19
C2324 vccd1.t72 vssa1 9.31e-19
C2325 vccd1.t69 vssa1 9.31e-19
C2326 vccd1.t62 vssa1 9.31e-19
C2327 vccd1.t42 vssa1 9.31e-19
C2328 vccd1.t71 vssa1 9.31e-19
C2329 vccd1.t53 vssa1 9.31e-19
C2330 vccd1.t57 vssa1 2.14e-19
C2331 vccd1.n72 vssa1 0.00144f
C2332 vccd1.n73 vssa1 7.34e-19
C2333 vccd1.n74 vssa1 0.00258f
C2334 vccd1.n75 vssa1 0.00132f
C2335 vccd1.t39 vssa1 1.9e-19
C2336 vccd1.t40 vssa1 1.9e-19
C2337 vccd1.n76 vssa1 4.7e-19
C2338 vccd1.t38 vssa1 0.00333f
C2339 vccd1.n77 vssa1 0.00179f
C2340 vccd1.n78 vssa1 4.7e-19
C2341 vccd1.n79 vssa1 3.38e-19
C2342 vccd1.n80 vssa1 1.04e-19
C2343 vccd1.n81 vssa1 3.42e-19
C2344 vccd1.t29 vssa1 1.9e-19
C2345 vccd1.t30 vssa1 1.9e-19
C2346 vccd1.n82 vssa1 4.7e-19
C2347 vccd1.t28 vssa1 0.00333f
C2348 vccd1.n83 vssa1 0.00179f
C2349 vccd1.n84 vssa1 4.7e-19
C2350 vccd1.n85 vssa1 7.2e-19
C2351 vccd1.n86 vssa1 0.00163f
C2352 vccd1.n87 vssa1 0.00154f
C2353 vccd1.n88 vssa1 0.00154f
C2354 vccd1.n89 vssa1 0.00154f
C2355 vccd1.n90 vssa1 0.00154f
C2356 vccd1.n91 vssa1 0.00154f
C2357 vccd1.n92 vssa1 0.00138f
C2358 vccd1.t3 vssa1 0.169f
C2359 vccd1.n93 vssa1 0.0498f
C2360 vccd1.n94 vssa1 3.3e-19
C2361 vccd1.n95 vssa1 0.00137f
C2362 vccd1.n96 vssa1 0.00154f
C2363 vccd1.n97 vssa1 0.00154f
C2364 vccd1.n98 vssa1 0.00154f
C2365 vccd1.n99 vssa1 0.00154f
C2366 vccd1.n100 vssa1 0.00154f
C2367 vccd1.n101 vssa1 0.00164f
C2368 vccd1.n102 vssa1 7.47e-19
C2369 vccd1.t5 vssa1 1.9e-19
C2370 vccd1.t4 vssa1 1.9e-19
C2371 vccd1.n103 vssa1 4.85e-19
C2372 vccd1.t2 vssa1 0.00333f
C2373 vccd1.n104 vssa1 0.00179f
C2374 vccd1.n105 vssa1 4.85e-19
C2375 vccd1.n106 vssa1 3.57e-19
C2376 vccd1.n107 vssa1 1.04e-19
C2377 vccd1.n108 vssa1 3.53e-19
C2378 vccd1.t27 vssa1 1.9e-19
C2379 vccd1.t26 vssa1 1.9e-19
C2380 vccd1.n109 vssa1 4.85e-19
C2381 vccd1.t24 vssa1 0.00333f
C2382 vccd1.n110 vssa1 0.00179f
C2383 vccd1.n111 vssa1 4.85e-19
C2384 vccd1.n112 vssa1 3.91e-19
C2385 vccd1.n113 vssa1 0.00138f
C2386 vccd1.n114 vssa1 7.46e-19
C2387 vccd1.t36 vssa1 4.27e-20
C2388 vccd1.n115 vssa1 5.47e-19
C2389 vccd1.n116 vssa1 0.00191f
C2390 vccd1.t35 vssa1 0.00134f
C2391 vccd1.n117 vssa1 0.00259f
C2392 vccd1.n118 vssa1 7.47e-19
C2393 vccd1.n119 vssa1 1.16e-19
C2394 vccd1.n120 vssa1 6.81e-19
C2395 vccd1.t18 vssa1 4.27e-20
C2396 vccd1.n121 vssa1 5.47e-19
C2397 vccd1.n122 vssa1 0.00191f
C2398 vccd1.t17 vssa1 0.00134f
C2399 vccd1.n123 vssa1 0.00259f
C2400 vccd1.n124 vssa1 0.0018f
C2401 vccd1.n125 vssa1 0.042f
C2402 vccd1.t7 vssa1 0.048f
C2403 vccd1.n126 vssa1 0.0399f
C2404 vccd1.n127 vssa1 0.00225f
C2405 vccd1.n128 vssa1 0.00174f
C2406 vccd1.t9 vssa1 4.27e-20
C2407 vccd1.n129 vssa1 5.47e-19
C2408 vccd1.n130 vssa1 0.00191f
C2409 vccd1.t6 vssa1 0.00134f
C2410 vccd1.n131 vssa1 0.0025f
C2411 vccd1.n132 vssa1 6.25e-19
C2412 vccd1.n133 vssa1 1.16e-19
C2413 vccd1.n134 vssa1 6.91e-19
C2414 vccd1.t23 vssa1 4.27e-20
C2415 vccd1.n135 vssa1 5.47e-19
C2416 vccd1.n136 vssa1 0.00191f
C2417 vccd1.t20 vssa1 0.00134f
C2418 vccd1.n137 vssa1 0.0025f
C2419 vccd1.n138 vssa1 0.00105f
C2420 vccd1.t63 vssa1 9.71e-19
C2421 vccd1.n139 vssa1 0.00166f
C2422 vccd1.t76 vssa1 9.71e-19
C2423 vccd1.n140 vssa1 0.00139f
C2424 vccd1.n141 vssa1 3.3e-19
C2425 vccd1.n142 vssa1 0.00278f
C2426 vccd1.n143 vssa1 0.0598f
C2427 vccd1.t25 vssa1 0.153f
C2428 vccd1.n144 vssa1 0.0505f
C2429 vccd1.n145 vssa1 0.0167f
C2430 vccd1.n146 vssa1 0.00957f
C2431 vccd1.n147 vssa1 2.47e-19
C2432 pmu_circuits_0.iref_2nA_0.iref_2nA_vref_0.DD vssa1 0.0057f
C2433 vccd1.n148 vssa1 0.00415f
C2434 vccd1.n149 vssa1 0.00805f
C2435 vccd1.n150 vssa1 0.0012f
C2436 vccd1.t55 vssa1 0.018f
C2437 vccd1.n151 vssa1 0.0176f
C2438 vccd1.t50 vssa1 0.018f
C2439 vccd1.n152 vssa1 0.0134f
C2440 vccd1.n153 vssa1 0.0014f
C2441 vccd1.n154 vssa1 0.00124f
C2442 vccd1.n155 vssa1 0.00123f
C2443 vccd1.n156 vssa1 7.62e-19
C2444 vccd1.n157 vssa1 0.00223f
C2445 vccd1.n159 vssa1 3.19e-19
C2446 vccd1.n160 vssa1 0.00139f
C2447 vccd1.n161 vssa1 0.0264f
C2448 pmu_circuits_0.iref_2nA_0.DD vssa1 0.252f
C2449 vccd1.n162 vssa1 0.272f
C2450 pmu_circuits_0.dd_01 vssa1 15.4f
C2451 a_337443_613718.n0 vssa1 1.26f
C2452 a_337443_613718.t3 vssa1 0.0123f
C2453 a_337443_613718.t4 vssa1 0.394f
C2454 a_337443_613718.t2 vssa1 0.394f
C2455 a_337443_613718.t1 vssa1 0.0122f
C2456 a_337443_613718.t5 vssa1 0.0122f
C2457 a_337443_613718.t0 vssa1 0.0122f
.ends


* NGSPICE file created from pmu_circuits.ext - technology: sky130A

.subckt pmu_circuits vref ldo_vs ldo_vb ldo_iref iref dd_02 ring_out ldo_out dd_01
+ ss
X0 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t5 iref_2nA_0.iref_2nA_igenerator_0.Vg ss.t126 ss.t125 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X1 dd_01.t20 a_1555_7968.t3 a_1555_7968.t4 dd_01.t18 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X2 dd_02.t36 ring_100mV_0.mdls_inv_2.IN a_7406_13329# ss.t192 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X3 ring_100mV_0.mdls_inv_5.OUT ring_100mV_0.mdls_inv_2.OUT a_9754_13622.t5 ss.t20 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X4 ss.t97 ldo_iref.t2 ldo_iref.t3 ss.t96 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X5 a_7406_11663# ring_100mV_0.mdls_inv_6.IN.t5 dd_02.t13 dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X6 dd_01.t31 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t3 a_1786_15962# dd_01.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X7 dd_01.t73 dd_01.t71 dd_01.t72 dd_01.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=2
X8 dd_01.t17 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t12 a_3482_12058# dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X9 dd_02.t40 ring_100mV_0.mdls_inv_3.OUT.t5 a_7406_14995# ss.t215 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X10 ss.t169 a_16150_16902.t6 vref.t3 ss.t168 sky130_fd_pr__nfet_01v8 ad=0.238 pd=2.22 as=0.238 ps=2.22 w=0.82 l=1.05
X11 ss.t24 ldo_iref.t4 a_14834_9380.t7 ss.t23 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X12 ring_100mV_0.mdls_inv_0.OUT.t3 ring_100mV_0.mdls_inv_0.IN a_9754_8624.t1 ss.t159 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X13 ring_100mV_0.mdls_inv_0.OUT.t2 ring_100mV_0.mdls_inv_0.IN a_9754_8624.t2 ss.t158 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X14 ring_100mV_0.mdls_inv_1.OUT.t2 ring_100mV_0.mdls_inv_0.OUT.t5 a_7406_8331# dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X15 dd_01.t32 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t4 a_1786_15962# dd_01.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X16 iref_2nA_0.iref_2nA_igenerator_0.VCTAT ss.t86 ss.t87 iref_2nA_0.iref_2nA_igenerator_0.VCTAT sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X17 dd_01.t75 a_15054_7578.t6 a_14490_9380.t1 dd_01.t74 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X18 ring_100mV_0.mdls_inv_1.OUT.t4 ring_100mV_0.mdls_inv_0.OUT.t6 a_5930_7513.t3 ss.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X19 ring_100mV_0.mdls_inv_1.OUT.t3 ring_100mV_0.mdls_inv_0.OUT.t7 a_5930_7513.t2 ss.t147 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X20 dd_01.t36 a_15054_7578.t2 a_15054_7578.t3 dd_01.t35 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X21 a_9754_11956.t6 ring_100mV_0.mdls_inv_5.OUT ss.t209 ss.t208 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X22 dd_01.t70 dd_01.t68 a_955_10311.t1 dd_01.t69 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X23 ring_out.t19 a_5712_16467.t10 ss.t7 ss.t6 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X24 a_5712_16467.t1 ring_100mV_0.mdls_inv_3.OUT.t6 dd_02.t42 dd_02.t41 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X25 iref_2nA_0.iref_2nA_igenerator_0.Vg a_n169_16287.t6 ss.t106 ss.t105 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X26 a_9754_14652# ring_100mV_0.mdls_inv_2.IN dd_02.t35 dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X27 dd_01.t67 dd_01.t64 dd_01.t66 dd_01.t65 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.258 ps=2.36 w=0.89 l=3.89
X28 a_9754_15288.t6 ring_100mV_0.mdls_inv_2.IN ss.t191 ss.t190 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X29 a_5930_7513.t5 ring_100mV_0.mdls_inv_0.OUT.t8 ss.t51 ss.t50 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X30 ss.t227 ring_100mV_0.mdls_inv_3.OUT.t7 a_5930_14177.t0 dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X31 a_5930_14177.t6 ring_100mV_0.mdls_inv_2.IN ss.t189 ss.t188 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X32 dd_02.t28 ring_100mV_0.mdls_inv_0.OUT.t9 a_9754_7988# ss.t146 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X33 dd_01.t63 dd_01.t61 dd_01.t62 dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=2
X34 ring_out.t18 a_5712_16467.t11 ss.t118 ss.t117 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X35 ring_100mV_0.mdls_inv_4.IN.t3 ring_100mV_0.mdls_inv_6.IN.t6 a_5930_10845.t2 ss.t130 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X36 dd_01.t38 a_14490_9380.t4 ldo_out.t4 dd_01.t37 sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.9 as=1.5 ps=10.9 w=5.17 l=0.37
X37 a_3482_8138.t9 a_n81_16487.t6 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t8 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X38 ring_100mV_0.mdls_inv_2.OUT ring_100mV_0.mdls_inv_2.IN a_9754_15288.t4 ss.t187 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X39 ss.t108 ring_100mV_0.mdls_inv_3.OUT.t8 a_5712_16467.t9 ss.t107 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X40 dd_01.t19 a_1555_7968.t1 a_1555_7968.t2 dd_01.t18 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X41 ring_100mV_0.mdls_inv_0.IN ring_100mV_0.mdls_inv_7.OUT a_9754_10290.t5 ss.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X42 ss.t144 ring_100mV_0.mdls_inv_0.OUT.t10 a_9754_8624.t0 dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X43 a_9754_13622.t1 ring_100mV_0.mdls_inv_2.OUT ss.t19 ss.t18 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X44 dd_01.t16 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t13 a_3482_8138.t19 dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X45 dd_01.t15 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t14 a_3482_12842# dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X46 ring_out.t17 a_5712_16467.t12 ss.t226 ss.t225 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X47 dd_02.t31 ring_100mV_0.mdls_inv_0.IN a_9754_9654# ss.t157 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X48 ring_100mV_0.mdls_inv_6.IN.t3 ring_100mV_0.mdls_inv_1.OUT.t5 a_5930_9179.t4 ss.t222 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X49 ss.t95 ss.t92 ss.t94 ss.t93 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=1.48 ps=10.8 w=5.1 l=0.66
X50 ss.t22 ring_100mV_0.mdls_inv_3.OUT.t9 a_5712_16467.t8 ss.t21 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X51 a_1786_16746# a_n81_16487.t7 iref_2nA_0.iref_2nA_igenerator_0.Vg dd_01.t24 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X52 w_583_11504# w_583_11504# ss.t8 w_583_11504# sky130_fd_pr__pfet_01v8_lvt ad=0.255 pd=2.34 as=0.255 ps=2.34 w=0.88 l=6.97
X53 ring_100mV_0.mdls_inv_2.IN ring_100mV_0.mdls_inv_4.IN.t5 a_7406_13329# dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X54 a_7406_8331# ring_100mV_0.mdls_inv_0.OUT.t11 dd_02.t43 dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X55 a_3482_8138.t8 a_n81_16487.t8 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t7 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X56 a_15054_7578.t5 ldo_iref.t5 ss.t41 ss.t40 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X57 iref_2nA_0.iref_2nA_igenerator_0.Vg a_n169_16287.t7 ss.t116 ss.t115 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X58 ss.t91 ss.t88 ss.t90 ss.t89 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0 ps=0 w=2.5 l=1
X59 dd_01.t14 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t15 a_3482_8138.t18 dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X60 dd_01.t21 a_16150_16902.t4 a_16150_16902.t5 ss.t47 sky130_fd_pr__nfet_01v8_lvt ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.89
X61 ring_100mV_0.mdls_inv_2.IN ring_100mV_0.mdls_inv_4.IN.t6 a_5930_12511.t5 ss.t171 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X62 a_3482_12842# a_n81_16487.t9 iref.t1 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X63 ring_100mV_0.mdls_inv_2.IN ring_100mV_0.mdls_inv_4.IN.t7 a_5930_12511.t4 ss.t148 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X64 dd_02.t11 ring_100mV_0.mdls_inv_4.IN.t8 a_7406_11663# ss.t37 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X65 dd_01.t13 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t16 a_3482_8138.t17 dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X66 dd_01.t28 a_16150_16902.t2 a_16150_16902.t3 ss.t109 sky130_fd_pr__nfet_01v8_lvt ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.89
X67 ring_100mV_0.mdls_inv_3.OUT.t3 ring_100mV_0.mdls_inv_2.IN a_7406_14995# dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X68 ss.t156 ring_100mV_0.mdls_inv_0.IN a_9754_10290.t6 dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X69 ring_100mV_0.mdls_inv_0.IN ring_100mV_0.mdls_inv_7.OUT a_9754_10290.t4 ss.t35 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X70 dd_02.t26 ring_100mV_0.mdls_inv_6.IN.t7 a_7406_9997# ss.t127 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X71 ring_out.t16 a_5712_16467.t13 ss.t100 ss.t99 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X72 a_9754_15288.t5 ring_100mV_0.mdls_inv_2.IN ss.t186 ss.t185 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X73 ring_out.t15 a_5712_16467.t14 ss.t104 ss.t103 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X74 ss.t207 ring_100mV_0.mdls_inv_5.OUT a_9754_13622.t6 dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X75 dd_02.t39 ring_100mV_0.mdls_inv_5.OUT a_9754_12986# ss.t206 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X76 dd_02.t23 a_5712_16467.t15 ring_out.t3 dd_02.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X77 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t4 iref_2nA_0.iref_2nA_igenerator_0.Vg ss.t124 ss.t123 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X78 ring_100mV_0.mdls_inv_0.OUT.t1 ring_100mV_0.mdls_inv_0.IN a_9754_8624.t6 ss.t155 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X79 dd_02.t7 ring_100mV_0.mdls_inv_2.OUT a_9754_14652# ss.t17 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X80 ring_100mV_0.mdls_inv_0.OUT.t0 ring_100mV_0.mdls_inv_0.IN a_9754_8624.t5 ss.t154 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X81 a_9754_11320# ring_100mV_0.mdls_inv_5.OUT dd_02.t38 dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X82 dd_01.t12 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t17 a_3482_8138.t16 dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X83 vref.t4 a_16150_16902.t0 a_16150_16902.t1 ss.t220 sky130_fd_pr__nfet_01v8_lvt ad=0.499 pd=4.02 as=0.499 ps=4.02 w=1.72 l=3.1
X84 vref.t2 vref.t0 vref.t1 dd_01.t76 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=8.6 ps=19.2 w=8.6 l=0.35
X85 ss.t85 ss.t82 ss.t84 ss.t83 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.725 ps=5.58 w=2.5 l=1
X86 a_9754_8624.t4 ring_100mV_0.mdls_inv_0.IN ss.t153 ss.t152 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X87 ring_100mV_0.mdls_inv_1.OUT.t1 ring_100mV_0.mdls_inv_0.OUT.t12 a_5930_7513.t1 ss.t161 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X88 ring_out.t14 a_5712_16467.t16 ss.t211 ss.t210 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X89 ring_100mV_0.mdls_inv_1.OUT.t0 ring_100mV_0.mdls_inv_0.OUT.t13 a_5930_7513.t0 ss.t160 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X90 a_3482_8138.t7 a_n81_16487.t10 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t1 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X91 a_1786_16746# a_n81_16487.t11 iref_2nA_0.iref_2nA_igenerator_0.Vg dd_01.t24 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X92 dd_01.t60 dd_01.t58 dd_01.t59 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=2
X93 a_3482_8138.t6 a_n81_16487.t12 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t10 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X94 a_7406_13329# ring_100mV_0.mdls_inv_4.IN.t9 dd_02.t14 dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X95 a_14834_9380.t1 ldo_vb.t0 a_14490_9380.t3 ss.t170 sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=5.19 l=1.43
X96 ring_100mV_0.mdls_inv_2.OUT ring_100mV_0.mdls_inv_2.IN a_9754_15288.t3 ss.t184 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X97 ring_100mV_0.mdls_inv_7.OUT ring_100mV_0.mdls_inv_5.OUT a_9754_11956.t4 ss.t205 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X98 ring_100mV_0.mdls_inv_2.OUT ring_100mV_0.mdls_inv_2.IN a_9754_15288.t2 ss.t183 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X99 ss.t102 ring_100mV_0.mdls_inv_4.IN.t10 a_5930_10845.t6 dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X100 ring_100mV_0.mdls_inv_0.OUT.t4 ring_100mV_0.mdls_inv_0.IN a_9754_7988# dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X101 ring_100mV_0.mdls_inv_0.IN ring_100mV_0.mdls_inv_7.OUT a_9754_10290.t3 ss.t34 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X102 ring_100mV_0.mdls_inv_3.OUT.t0 ring_100mV_0.mdls_inv_2.IN a_5930_14177.t4 ss.t182 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X103 ring_100mV_0.mdls_inv_0.IN ring_100mV_0.mdls_inv_7.OUT a_9754_10290.t2 ss.t33 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X104 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t1 iref_2nA_0.iref_2nA_igenerator_0.Vg a_828_14113# ss.t122 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X105 ss.t57 ldo_iref.t6 a_14834_9380.t6 ss.t56 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X106 dd_02.t12 ring_100mV_0.mdls_inv_4.IN.t11 a_7406_11663# ss.t44 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X107 ss.t16 ring_100mV_0.mdls_inv_2.OUT a_9754_15288.t0 dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X108 ring_100mV_0.mdls_inv_6.IN.t0 ring_100mV_0.mdls_inv_1.OUT.t6 a_7406_9997# dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X109 ring_100mV_0.mdls_inv_6.IN.t1 ring_100mV_0.mdls_inv_1.OUT.t7 a_5930_9179.t3 ss.t112 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X110 ring_100mV_0.mdls_inv_6.IN.t2 ring_100mV_0.mdls_inv_1.OUT.t8 a_5930_9179.t2 ss.t214 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X111 ring_100mV_0.mdls_inv_2.OUT ring_100mV_0.mdls_inv_2.IN a_9754_15288.t1 ss.t181 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X112 a_n169_16287.t4 a_n169_16287.t3 ss.t120 ss.t119 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X113 dd_02.t3 ring_100mV_0.mdls_inv_3.OUT.t10 a_7406_14995# ss.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X114 ss.t139 ldo_iref.t7 a_15054_7578.t4 ss.t138 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X115 dd_01.t11 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t18 a_3482_8138.t15 dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X116 ring_out.t13 a_5712_16467.t17 ss.t198 ss.t197 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X117 dd_02.t1 ring_100mV_0.mdls_inv_3.OUT.t11 a_5712_16467.t0 dd_02.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X118 a_828_14113# iref_2nA_0.iref_2nA_igenerator_0.VCTAT ss.t63 ss.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=5
X119 dd_02.t27 ring_100mV_0.mdls_inv_1.OUT.t9 a_7406_8331# ss.t145 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X120 dd_01.t25 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t5 a_1786_16746# dd_01.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X121 a_3482_8138.t5 a_n81_16487.t13 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t3 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X122 a_3482_12058# a_n81_16487.t14 a_n169_16287.t0 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X123 a_955_10311.t0 w_583_11504# iref_2nA_0.iref_2nA_igenerator_0.VCTAT dd_01.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.995 pd=7.44 as=0.995 ps=7.44 w=3.43 l=2.77
X124 ss.t5 ring_100mV_0.mdls_inv_3.OUT.t12 a_5712_16467.t7 ss.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X125 dd_01.t57 dd_01.t54 dd_01.t56 dd_01.t55 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0 ps=0 w=0.89 l=3.89
X126 a_3482_8138.t4 a_n81_16487.t15 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t6 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X127 a_5930_12511.t1 ring_100mV_0.mdls_inv_4.IN.t12 ss.t134 ss.t133 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X128 dd_01.t27 a_15054_7578.t0 a_15054_7578.t1 dd_01.t26 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X129 ring_100mV_0.mdls_inv_5.OUT ring_100mV_0.mdls_inv_2.OUT a_9754_12986# dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X130 a_5930_9179.t6 ring_100mV_0.mdls_inv_1.OUT.t10 ss.t59 ss.t58 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X131 ring_100mV_0.mdls_inv_6.IN.t4 ring_100mV_0.mdls_inv_1.OUT.t11 a_5930_9179.t1 ss.t232 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X132 dd_01.t30 a_15054_7578.t7 a_14490_9380.t0 dd_01.t29 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X133 a_n81_16487.t5 a_n169_16287.t8 ss.t213 ss.t212 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X134 dd_02.t10 ring_100mV_0.mdls_inv_7.OUT a_9754_11320# ss.t32 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X135 dd_01.t53 dd_01.t51 dd_01.t52 dd_01.t24 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=2
X136 a_9754_7988# ring_100mV_0.mdls_inv_0.IN dd_02.t30 dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X137 ring_100mV_0.mdls_inv_4.IN.t4 ring_100mV_0.mdls_inv_6.IN.t8 a_7406_11663# dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X138 ss.t81 ss.t78 ss.t80 ss.t79 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0 ps=0 w=2.5 l=1
X139 ring_out.t12 a_5712_16467.t18 ss.t46 ss.t45 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X140 dd_01.t10 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t19 a_3482_8138.t14 dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X141 ring_out.t2 a_5712_16467.t19 dd_02.t17 dd_02.t16 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X142 dd_02.t29 ring_100mV_0.mdls_inv_0.IN a_9754_9654# ss.t151 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X143 ring_100mV_0.mdls_inv_2.OUT ring_100mV_0.mdls_inv_2.IN a_9754_14652# dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X144 a_14834_9380.t5 ldo_iref.t8 ss.t141 ss.t140 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X145 a_14834_9380.t0 ldo_vb.t1 a_14490_9380.t2 ss.t170 sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=5.19 l=1.43
X146 a_5930_10845.t4 ring_100mV_0.mdls_inv_6.IN.t9 ss.t194 ss.t193 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X147 a_5930_7513.t4 ring_100mV_0.mdls_inv_0.OUT.t14 ss.t196 ss.t195 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X148 dd_01.t23 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t6 a_1786_16746# dd_01.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X149 ring_out.t11 a_5712_16467.t20 ss.t53 ss.t52 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X150 dd_02.t34 ring_100mV_0.mdls_inv_2.IN a_7406_13329# ss.t180 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X151 a_14834_9380.t4 ldo_iref.t9 ss.t219 ss.t218 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X152 dd_01.t34 a_955_10311.t2 w_583_11504# dd_01.t33 sky130_fd_pr__pfet_01v8 ad=0.687 pd=5.32 as=0.687 ps=5.32 w=2.37 l=4.38
X153 dd_01.t9 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t20 a_3482_12842# dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X154 ring_100mV_0.mdls_inv_3.OUT.t2 ring_100mV_0.mdls_inv_2.IN a_5930_14177.t3 ss.t179 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X155 a_7406_9997# ring_100mV_0.mdls_inv_1.OUT.t12 dd_02.t15 dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X156 ring_100mV_0.mdls_inv_4.IN.t2 ring_100mV_0.mdls_inv_6.IN.t10 a_5930_10845.t5 ss.t135 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X157 ss.t39 ring_100mV_0.mdls_inv_3.OUT.t13 a_5712_16467.t6 ss.t38 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X158 ring_100mV_0.mdls_inv_3.OUT.t4 ring_100mV_0.mdls_inv_2.IN a_5930_14177.t2 ss.t178 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X159 a_n169_16287.t2 a_n169_16287.t1 ss.t55 ss.t54 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X160 ring_100mV_0.mdls_inv_7.OUT ring_100mV_0.mdls_inv_5.OUT a_9754_11956.t3 ss.t204 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X161 dd_01.t50 dd_01.t48 dd_01.t49 dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=2
X162 ring_out.t10 a_5712_16467.t21 ss.t167 ss.t166 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X163 ring_100mV_0.mdls_inv_7.OUT ring_100mV_0.mdls_inv_5.OUT a_9754_11956.t2 ss.t203 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X164 a_3482_12058# a_n81_16487.t16 a_n169_16287.t5 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X165 ring_100mV_0.mdls_inv_3.OUT.t1 ring_100mV_0.mdls_inv_2.IN a_5930_14177.t1 ss.t177 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X166 ss.t129 ring_100mV_0.mdls_inv_3.OUT.t14 a_5712_16467.t5 ss.t128 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X167 a_9754_12986# ring_100mV_0.mdls_inv_2.OUT dd_02.t6 dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X168 a_9754_13622.t0 ring_100mV_0.mdls_inv_2.OUT ss.t15 ss.t14 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X169 ss.t31 ring_100mV_0.mdls_inv_7.OUT a_9754_11956.t0 dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X170 dd_02.t9 ring_100mV_0.mdls_inv_7.OUT a_9754_11320# ss.t30 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X171 a_1555_7968.t5 a_n81_16487.t2 a_n81_16487.t3 dd_01.t1 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X172 a_5930_9179.t5 ring_100mV_0.mdls_inv_1.OUT.t13 ss.t111 ss.t110 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X173 dd_01.t8 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t21 a_3482_8138.t13 dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X174 ring_out.t9 a_5712_16467.t22 ss.t132 ss.t131 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X175 dd_02.t4 ring_100mV_0.mdls_inv_2.OUT a_9754_14652# ss.t13 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X176 dd_01.t7 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t22 a_3482_8138.t12 dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X177 dd_02.t18 ring_100mV_0.mdls_inv_0.OUT.t15 a_9754_7988# ss.t61 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X178 ring_100mV_0.mdls_inv_5.OUT ring_100mV_0.mdls_inv_2.OUT a_9754_13622.t4 ss.t12 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X179 iref_2nA_0.iref_2nA_igenerator_0.VCTAT ss.t70 ss.t71 iref_2nA_0.iref_2nA_igenerator_0.VCTAT sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X180 ring_100mV_0.mdls_inv_5.OUT ring_100mV_0.mdls_inv_2.OUT a_9754_13622.t3 ss.t11 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X181 a_9754_10290.t1 ring_100mV_0.mdls_inv_7.OUT ss.t29 ss.t28 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X182 ring_100mV_0.mdls_inv_0.IN ring_100mV_0.mdls_inv_7.OUT a_9754_9654# dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X183 a_9754_11956.t5 ring_100mV_0.mdls_inv_5.OUT ss.t202 ss.t201 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X184 a_1786_15962# a_n81_16487.t17 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t2 dd_01.t24 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X185 a_n81_16487.t4 a_n169_16287.t9 ss.t2 ss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X186 dd_01.t47 dd_01.t45 dd_01.t46 dd_01.t24 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=2
X187 dd_01.t44 dd_01.t42 dd_01.t43 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=2
X188 ring_out.t8 a_5712_16467.t23 ss.t231 ss.t230 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X189 iref_2nA_0.iref_2nA_igenerator_0.VCTAT ss.t76 ss.t77 iref_2nA_0.iref_2nA_igenerator_0.VCTAT sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X190 dd_02.t25 a_5712_16467.t24 ring_out.t1 dd_02.t24 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X191 ldo_out.t2 ldo_vs.t0 a_14834_9380.t3 ldo_out.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.76 pd=12.7 as=1.76 ps=12.7 w=6.07 l=1.27
X192 a_7406_14995# ring_100mV_0.mdls_inv_2.IN dd_02.t33 dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X193 dd_01.t6 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t23 a_3482_8138.t11 dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X194 ss.t163 ring_100mV_0.mdls_inv_3.OUT.t15 a_5712_16467.t4 ss.t162 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X195 dd_01.t41 dd_01.t39 dd_01.t40 dd_01.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=2
X196 a_1786_15962# a_n81_16487.t18 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t0 dd_01.t24 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X197 ss.t75 ss.t72 ss.t74 ss.t73 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=0 ps=0 w=5.1 l=0.66
X198 a_3482_8138.t3 a_n81_16487.t19 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t9 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X199 a_3482_12842# a_n81_16487.t20 iref.t0 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X200 dd_01.t5 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t24 a_3482_8138.t10 dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X201 dd_01.t4 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t25 a_3482_12058# dd_01.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X202 ring_out.t7 a_5712_16467.t25 ss.t217 ss.t216 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X203 a_9754_8624.t3 ring_100mV_0.mdls_inv_0.IN ss.t150 ss.t149 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X204 ss.t221 ring_100mV_0.mdls_inv_1.OUT.t14 a_5930_7513.t6 dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X205 ss.t173 ring_100mV_0.mdls_inv_3.OUT.t16 a_5712_16467.t3 ss.t172 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X206 a_14490_9380.t5 ldo_out.t3 sky130_fd_pr__cap_mim_m3_1 l=15 w=4
X207 dd_02.t19 ring_100mV_0.mdls_inv_1.OUT.t15 a_7406_8331# ss.t98 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X208 a_1555_7968.t0 a_n81_16487.t0 a_n81_16487.t1 dd_01.t1 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X209 ring_100mV_0.mdls_inv_7.OUT ring_100mV_0.mdls_inv_5.OUT a_9754_11320# dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X210 ring_100mV_0.mdls_inv_7.OUT ring_100mV_0.mdls_inv_5.OUT a_9754_11956.t1 ss.t200 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X211 dd_02.t32 ring_100mV_0.mdls_inv_6.IN.t11 a_7406_9997# ss.t165 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X212 ring_100mV_0.mdls_inv_4.IN.t1 ring_100mV_0.mdls_inv_6.IN.t12 a_5930_10845.t1 ss.t25 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X213 a_3482_8138.t2 a_n81_16487.t21 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t11 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X214 dd_02.t37 ring_100mV_0.mdls_inv_5.OUT a_9754_12986# ss.t199 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
X215 a_5930_10845.t3 ring_100mV_0.mdls_inv_6.IN.t13 ss.t49 ss.t48 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X216 ring_100mV_0.mdls_inv_4.IN.t0 ring_100mV_0.mdls_inv_6.IN.t14 a_5930_10845.t0 ss.t60 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X217 iref_2nA_0.iref_2nA_igenerator_0.Ip1 iref_2nA_0.iref_2nA_igenerator_0.Vg a_828_14113# ss.t121 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X218 ring_out.t6 a_5712_16467.t26 ss.t224 ss.t223 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X219 ring_out.t5 a_5712_16467.t27 ss.t229 ss.t228 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X220 a_5930_14177.t5 ring_100mV_0.mdls_inv_2.IN ss.t176 ss.t175 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X221 ldo_out.t1 ldo_vs.t1 a_14834_9380.t2 ldo_out.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.76 pd=12.7 as=1.76 ps=12.7 w=6.07 l=1.27
X222 ring_out.t0 a_5712_16467.t28 dd_02.t21 dd_02.t20 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X223 a_3482_8138.t1 a_n81_16487.t22 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t2 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X224 a_9754_10290.t0 ring_100mV_0.mdls_inv_7.OUT ss.t27 ss.t26 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X225 a_3482_8138.t0 a_n81_16487.t23 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t0 dd_01.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
X226 ss.t3 ring_100mV_0.mdls_inv_6.IN.t15 a_5930_9179.t0 dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X227 a_9754_9654# ring_100mV_0.mdls_inv_7.OUT dd_02.t8 dd_02.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X228 iref_2nA_0.iref_2nA_igenerator_0.VCTAT ss.t68 ss.t69 iref_2nA_0.iref_2nA_igenerator_0.VCTAT sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X229 ring_out.t4 a_5712_16467.t29 ss.t114 ss.t113 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X230 ring_100mV_0.mdls_inv_2.IN ring_100mV_0.mdls_inv_4.IN.t13 a_5930_12511.t3 ss.t164 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X231 ring_100mV_0.mdls_inv_2.IN ring_100mV_0.mdls_inv_4.IN.t14 a_5930_12511.t2 ss.t101 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X232 ss.t174 ring_100mV_0.mdls_inv_2.IN a_5930_12511.t6 dd_02.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
X233 ldo_iref.t1 ldo_iref.t0 ss.t143 ss.t142 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X234 ss.t67 ss.t64 ss.t66 ss.t65 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.725 ps=5.58 w=2.5 l=1
X235 ss.t137 ring_100mV_0.mdls_inv_3.OUT.t17 a_5712_16467.t2 ss.t136 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
X236 a_5930_12511.t0 ring_100mV_0.mdls_inv_4.IN.t15 ss.t43 ss.t42 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
X237 ring_100mV_0.mdls_inv_5.OUT ring_100mV_0.mdls_inv_2.OUT a_9754_13622.t2 ss.t10 sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
R0 ss.n223 ss.n222 13074
R1 ss.n427 ss.n426 8070.56
R2 ss.n308 ss.n307 5645.54
R3 ss.n433 ss.n432 5504.01
R4 ss.n375 ss.n374 2131.18
R5 ss.n377 ss.n376 2131.18
R6 ss.n259 ss.n258 2131.18
R7 ss.n261 ss.n260 2131.18
R8 ss.n333 ss.n330 1772.94
R9 ss.n221 ss.n218 1549.06
R10 ss.n427 ss.n425 1421.99
R11 ss.n103 ss.n102 1332.51
R12 ss.n287 ss.n274 1303.68
R13 ss.n421 ss.n375 1093.73
R14 ss.n365 ss.n259 1093.73
R15 ss.n255 ss.n254 1050.42
R16 ss.n9 ss.n7 1039.43
R17 ss.n421 ss.n377 1037.45
R18 ss.n365 ss.n261 1037.45
R19 ss.n113 ss.n112 1022.2
R20 ss.n211 ss.n209 892.788
R21 ss.t79 ss.t1 873.699
R22 ss.t119 ss.t115 873.699
R23 ss.t54 ss.t105 873.699
R24 ss.t65 ss.t212 873.699
R25 ss.n339 ss.n294 770.619
R26 ss.n393 ss.n392 691.729
R27 ss.n32 ss.t65 657.375
R28 ss.n317 ss.n315 604.529
R29 ss.n50 ss.t79 569.165
R30 ss.t6 ss.t131 568.843
R31 ss.t197 ss.t223 568.843
R32 ss.t223 ss.t99 568.843
R33 ss.t228 ss.t45 568.843
R34 ss.t103 ss.t228 568.843
R35 ss.n366 ss.n365 547.604
R36 ss.n220 ss.n219 515.481
R37 ss.t73 ss.t138 482.06
R38 ss.t23 ss.t56 482.06
R39 ss.n44 ss.t119 464.154
R40 ss.n126 ss.t168 433.62
R41 ss.n423 ss.n422 408.563
R42 ss.n280 ss.n277 404.93
R43 ss.n214 ss.n213 400.829
R44 ss.n28 ss.t122 367.111
R45 ss.n43 ss.t54 352.841
R46 ss.t42 ss.t164 346.818
R47 ss.t60 ss.t193 346.818
R48 ss.t195 ss.t0 346.818
R49 ss.n137 ss.n101 344
R50 ss.n129 ss.t47 342.469
R51 ss.t183 ss.t185 338.611
R52 ss.t12 ss.t18 338.611
R53 ss.t159 ss.t149 338.611
R54 ss.n136 ss.n105 333.382
R55 ss.n316 ss.t73 309.724
R56 ss.t62 ss.t121 306.812
R57 ss.t9 ss.t215 296.988
R58 ss.t37 ss.t44 296.988
R59 ss.t127 ss.t165 296.988
R60 ss.t145 ss.t98 296.988
R61 ss.t13 ss.t17 289.961
R62 ss.t199 ss.t206 289.961
R63 ss.n256 ss.t51 285.935
R64 ss.n248 ss.t59 285.935
R65 ss.n418 ss.t49 285.935
R66 ss.n397 ss.t134 285.935
R67 ss.n384 ss.t176 285.935
R68 ss.n85 ss.t191 285.935
R69 ss.n264 ss.t15 285.935
R70 ss.n362 ss.t209 285.935
R71 ss.n342 ss.t29 285.935
R72 ss.n257 ss.t153 285.935
R73 ss.n138 ss.t6 285.844
R74 ss.t179 ss.t175 283.036
R75 ss.t133 ss.t148 283.036
R76 ss.t214 ss.t58 283.036
R77 ss.t50 ss.t160 283.036
R78 ss.n138 ss.t197 283
R79 ss.t184 ss.t190 276.339
R80 ss.t14 ss.t20 276.339
R81 ss.n311 ss.n310 264.834
R82 ss.n395 ss.t192 256.127
R83 ss.t142 ss.t218 253.639
R84 ss.t40 ss.t140 253.639
R85 ss.n332 ss.t154 252.986
R86 ss.t162 ss.t117 243.62
R87 ss.t107 ss.t52 243.62
R88 ss.n166 ss.t177 238.189
R89 ss.t171 ss.n389 238.189
R90 ss.t130 ss.n407 238.189
R91 ss.n412 ss.t232 238.189
R92 ss.t161 ss.n253 238.189
R93 ss.n201 ss.n200 234.1
R94 ss.n88 ss.t181 232.553
R95 ss.t200 ss.n273 232.553
R96 ss.n135 ss.n108 226.969
R97 ss.n295 ss.t94 224.56
R98 ss.n288 ss.t30 221.85
R99 ss.n312 ss.t75 220.899
R100 ss.n298 ss.t23 218.132
R101 ss.n183 ss.n182 216.345
R102 ss.n420 ss.t25 214.27
R103 ss.n30 ss.n17 214.236
R104 ss.n352 ss.t155 214.065
R105 ss.n364 ss.t204 209.2
R106 ss.n22 ss.n20 207.369
R107 ss.n295 ss.t92 206.381
R108 ss.n321 ss.t72 206.317
R109 ss.n126 ss.t109 203.137
R110 ss.n176 ss.n70 200.833
R111 ss.n156 ss.t136 192.102
R112 ss.n285 ss.n280 192
R113 ss.t203 ss.t170 182.929
R114 ss.n26 ss.n25 179.953
R115 ss.n285 ss.n284 169.912
R116 ss.n182 ss.n179 163.743
R117 ss.n143 ss.t103 163.542
R118 ss.n292 ss.n291 162.329
R119 ss.n135 ss.n128 161.262
R120 ss.t21 ss.n175 160.667
R121 ss.t170 ss.t201 155.684
R122 ss.n148 ss.n147 148.107
R123 ss.t170 ss.t28 142.061
R124 ss.n301 ss.t142 142.038
R125 ss.n431 ss.n241 139.751
R126 ss.n87 ss.n86 139.143
R127 ss.t96 ss.n298 138.868
R128 ss.n208 ss.t124 135.946
R129 ss.n25 ss.t126 135.635
R130 ss.t170 ss.t34 134.278
R131 ss.n100 ss.n96 133.885
R132 ss.n439 ss.n183 132.236
R133 ss.n237 ss.t70 128.282
R134 ss.n306 ss.t139 127.653
R135 ss.n305 ss.t57 127.653
R136 ss.n296 ss.t24 127.653
R137 ss.n297 ss.t97 127.653
R138 ss.n304 ss.t143 127.653
R139 ss.n325 ss.t219 127.653
R140 ss.n326 ss.t141 127.653
R141 ss.n327 ss.t41 127.653
R142 ss.n227 ss.t68 127.34
R143 ss.n234 ss.t86 127.338
R144 ss.n282 ss.t35 126.493
R145 ss.n147 ss.n100 120.156
R146 ss.n2 ss.n1 118.558
R147 ss.n197 ss.n196 118.558
R148 ss.n249 ss.n248 113.725
R149 ss.n418 ss.n417 113.725
R150 ss.n398 ss.n397 113.725
R151 ss.n385 ss.n384 113.725
R152 ss.n85 ss.n84 113.725
R153 ss.n268 ss.n264 113.725
R154 ss.n362 ss.n361 113.725
R155 ss.n346 ss.n342 113.725
R156 ss.n210 ss.t83 113.504
R157 ss.n241 ss.n238 113.139
R158 ss.n322 ss.n306 112.356
R159 ss.n301 ss.t96 111.602
R160 ss.n198 ss.n195 110.448
R161 ss.n189 ss.n184 109.371
R162 ss.n46 ss.n36 108.484
R163 ss.n47 ss.n46 107.469
R164 ss.n282 ss.n281 106.059
R165 ss.t117 ss.t107 105.656
R166 ss.t52 ss.t38 105.656
R167 ss.t136 ss.t113 105.656
R168 ss.t210 ss.t4 105.656
R169 ss.t172 ss.t216 105.656
R170 ss.t225 ss.t21 105.656
R171 ss.t166 ss.t128 105.656
R172 ss.n431 ss.n430 102.694
R173 ss.n136 ss.n135 101.73
R174 ss.n218 ss.n215 99.3424
R175 ss.n73 ring_100mV_0.mdls_inv_2.SS 98.1054
R176 ss.n184 ss.t2 96.1374
R177 ss.n37 ss.t116 96.1374
R178 ss.n38 ss.t120 96.1374
R179 ss.n40 ss.t55 96.1374
R180 ss.n39 ss.t106 96.1374
R181 ss.n193 ss.t213 96.1374
R182 ss.n204 ss.t123 95.7683
R183 ss.n49 ss.n48 95.624
R184 ss.n392 ss.n47 95.2868
R185 ss.n194 ss.n193 92.7541
R186 ss.n383 ss.t182 84.7117
R187 ss.n396 ss.t101 84.7117
R188 ss.t135 ss.n419 84.7117
R189 ss.n247 ss.t222 84.7117
R190 ss.n255 ss.t147 84.7117
R191 ss.n286 ss.n285 84.7064
R192 ss.n368 ss.n257 83.6449
R193 ss.n372 ss.n256 83.6449
R194 ss.n175 ss.t166 82.9535
R195 ss.t187 ss.n87 82.7073
R196 ss.t205 ss.n363 82.7073
R197 ss.n341 ss.t36 82.7073
R198 ss.t158 ss.n331 82.7073
R199 ss.n424 ss.n423 82.5178
R200 ss.n38 ss.n37 77.1715
R201 ss.n40 ss.n39 77.1715
R202 ss.n123 ss.n122 76.2307
R203 ss.t175 ss.t178 75.7423
R204 ss.t164 ss.t133 75.7423
R205 ss.t48 ss.t60 75.7423
R206 ss.t58 ss.t112 75.7423
R207 ss.t0 ss.t50 75.7423
R208 ss.n24 ss.n23 75.2946
R209 ss.t190 ss.t183 73.9501
R210 ss.t208 ss.t203 73.9501
R211 ss.t28 ss.t33 73.9501
R212 ss.t152 ss.t159 73.9501
R213 ss.n2 ss.t64 73.5085
R214 ss.n197 ss.t82 73.5085
R215 ss.n5 ss.t88 73.5085
R216 ss.n185 ss.t78 73.5085
R217 ss.n5 ss.n4 73.2527
R218 ss.n186 ss.n185 73.2527
R219 ss.n31 ss.n30 72.0663
R220 ss.n438 ss.n437 68.8161
R221 ss.n420 ss.t48 68.7661
R222 ss.t32 ss.n288 68.112
R223 ss.n364 ss.t208 67.1389
R224 ss.n207 ss.n206 67.0123
R225 ss.n198 ss.n197 65.2057
R226 ss.n228 ss.t76 64.4538
R227 ss.n28 ss.t62 63.8457
R228 ss.n324 ss.n323 62.5845
R229 ss.n41 ss.n40 61.5889
R230 ss.n67 ss.t230 61.1237
R231 ss.n306 ss.n305 60.9529
R232 ss.n297 ss.n296 60.9529
R233 ss.t215 ss.t179 57.8034
R234 ss.t148 ss.t180 57.8034
R235 ss.t25 ss.t37 57.8034
R236 ss.t165 ss.t214 57.8034
R237 ss.t160 ss.t145 57.8034
R238 ss.n44 ss.n43 56.7069
R239 ss.t17 ss.t184 56.4357
R240 ss.t20 ss.t199 56.4357
R241 ss.t204 ss.t32 56.4357
R242 ss.t34 ss.t157 56.4357
R243 ss.t154 ss.t61 56.4357
R244 ss.n278 ss.t14 55.4627
R245 ring_100mV_0.mdls_inv_5.SS ss.n82 55.2813
R246 ring_100mV_0.mdls_inv_7.SS ss.n266 55.2813
R247 ring_100mV_0.mdls_inv_9.SS ss.n359 55.2813
R248 ring_100mV_0.mdls_inv_0.SS ss.n344 55.2813
R249 ss.n304 ss.n303 54.7053
R250 ss.n156 ss.t210 51.5187
R251 ring_100mV_0.mdls_inv_1.SS ss.n245 51.4565
R252 ss.n409 ring_100mV_0.mdls_inv_8.SS 51.4565
R253 ss.n400 ring_100mV_0.mdls_inv_6.SS 51.4565
R254 ring_100mV_0.mdls_inv_4.SS ss.n381 51.4565
R255 ss.n303 ss.n297 47.2386
R256 iref_2nA_0.iref_2nA_vref_0.SS ss.n224 47.1531
R257 ss.n3 ss.n0 47.1193
R258 ss.n187 ss.n186 47.1193
R259 ss.n436 ss.n212 46.7366
R260 ss.n225 iref_2nA_0.iref_2nA_vref_0.SS 45.8398
R261 ss.n25 ss.n24 45.4822
R262 ss.n94 ring_100mV_0.mdls_inv_2.SS 45.3694
R263 ss.n159 ss.n70 44.5387
R264 ss.n67 ss.t162 44.5331
R265 ss.n165 ss.n163 43.7783
R266 ss.n212 ss.n208 43.4171
R267 ss.n124 ss.n123 42.7248
R268 ss.n329 ss.n328 42.0106
R269 ss.n74 ss.n72 41.5894
R270 ss.t180 ss.n395 40.8612
R271 ss.n335 ss.n334 40.2265
R272 ss.n8 ss.t89 39.017
R273 ss.n84 ss.n75 38.6565
R274 ss.n269 ss.n268 38.6565
R275 ss.n361 ss.n353 38.6565
R276 ss.n347 ss.n346 38.6565
R277 ss.n250 ss.n249 38.5285
R278 ss.n417 ss.n416 38.5285
R279 ss.n386 ss.n385 38.5285
R280 ss.n167 ss.n166 37.8714
R281 ss.n389 ss.n388 37.8714
R282 ss.n407 ss.n406 37.8714
R283 ss.n414 ss.n412 37.8714
R284 ss.n253 ss.n252 37.8714
R285 ss.n12 ss.n11 37.8672
R286 ss.n12 ss.n10 37.109
R287 ss.n89 ss.n88 36.9753
R288 ss.n79 ss.n77 36.9753
R289 ss.n273 ss.n272 36.9753
R290 ss.n351 ss.n350 36.9753
R291 ss.n435 ss.n431 34.3363
R292 ss.n141 ss.n140 34.3018
R293 ss.n178 ss.n69 33.7524
R294 ss.n230 ss.t8 33.5458
R295 ss.n430 ss.n429 33.4393
R296 ss.n321 ss.n320 31.5524
R297 ss.n224 ss.n223 30.8191
R298 ss.n173 ss.n172 30.1042
R299 ss.n73 ss.t16 29.6448
R300 ss.n75 ss.t207 29.6448
R301 ss.n269 ss.t31 29.6448
R302 ss.n353 ss.t156 29.6448
R303 ss.n347 ss.t144 29.6448
R304 ss.n250 ss.t221 29.6447
R305 ss.n416 ss.t3 29.6447
R306 ss.n404 ss.t102 29.6447
R307 ss.n386 ss.t174 29.6447
R308 ss.n164 ss.t227 29.6447
R309 ss.n318 ss.n314 29.615
R310 ss.n423 ss.n373 29.0262
R311 ss.n70 ss.t172 28.8157
R312 ss.n437 ss.n436 28.8057
R313 ss.n21 ss.t125 28.3762
R314 ss.n324 ss.n304 28.191
R315 ss.n208 ss.n207 27.9094
R316 ss ss.t63 27.542
R317 vref01_0.SS ss.t169 26.8053
R318 ss.n336 ss.n335 26.5148
R319 ss.n225 ss.n217 26.1475
R320 ss.n3 ss.n2 26.1338
R321 ss.n191 ss.n190 26.1338
R322 ss.n35 ss.n31 24.043
R323 ss.n249 ss.n246 23.5607
R324 ss.n417 ss.n408 23.5607
R325 ss.n399 ss.n398 23.5607
R326 ss.n385 ss.n382 23.5607
R327 ss.n84 ss.n83 23.5607
R328 ss.n268 ss.n267 23.5607
R329 ss.n361 ss.n360 23.5607
R330 ss.n346 ss.n345 23.5607
R331 ss.t168 ss.t220 23.4394
R332 ss.n145 ss.n144 23.2318
R333 ss.n185 ss.n49 22.9338
R334 ss.n332 ss.t93 22.38
R335 ss.n36 ss.n3 21.6894
R336 ss.n338 ss.n337 20.3299
R337 ss.n17 ss.n5 19.9116
R338 ss.n140 ss.n137 18.8176
R339 ss.n98 ss.n97 18.4879
R340 ss.n278 ss.t12 18.4879
R341 ss.n352 ss.n351 18.4879
R342 ss.n436 ss.n435 18.2892
R343 ss.n7 ss.n6 18.1452
R344 ss.n192 ss.n191 17.9561
R345 ss.n372 ss.n371 17.6946
R346 ss.n441 ss.n49 17.4227
R347 ss.n144 ss.n143 17.0658
R348 ss.n371 ss.n368 16.2044
R349 ss.n13 ss.n12 16.0163
R350 ss.n35 ss.n34 16.0005
R351 ss.n41 ss.n38 15.5831
R352 ss.n367 ss.n366 15.3949
R353 ss.n229 ss.t77 14.906
R354 ss.n236 ss.t71 14.7432
R355 ss.n233 ss.t87 14.7432
R356 ss.n231 ss.t69 14.7432
R357 ss.n96 ss.n95 14.6846
R358 ss.t170 ss.n352 14.5847
R359 ss.n176 ss.t225 13.9715
R360 ss.n17 ss.n16 13.9355
R361 ss.n335 ss.n295 13.0318
R362 ss.n438 ss.n189 12.8666
R363 ss.n170 ss.n169 12.6654
R364 ss.n437 ss.n194 12.5496
R365 ss.t182 ss.t188 11.9597
R366 ss.t101 ss.t42 11.9597
R367 ss.t193 ss.t135 11.9597
R368 ss.t222 ss.t110 11.9597
R369 ss.t147 ss.t195 11.9597
R370 ss.t185 ss.t187 11.6767
R371 ss.t18 ss.t11 11.6767
R372 ss.t201 ss.t205 11.6767
R373 ss.t36 ss.t26 11.6767
R374 ss.t149 ss.t158 11.6767
R375 ss.n171 ring_100mV_0.ring_100mV_buffer_0.SS 11.5307
R376 ss.n179 ring_100mV_0.ring_100mV_buffer_0.SS 10.1931
R377 ss.n158 ring_100mV_0.mdls_inv_3.SS 10.059
R378 ss.n439 ss.n438 9.47205
R379 ss.n123 vref01_0.SS 9.30283
R380 ss.n117 ss.n111 9.1686
R381 ss.n246 ring_100mV_0.mdls_inv_1.SS 8.9248
R382 ring_100mV_0.mdls_inv_8.SS ss.n408 8.9248
R383 ring_100mV_0.mdls_inv_6.SS ss.n399 8.9248
R384 ss.n382 ring_100mV_0.mdls_inv_4.SS 8.9248
R385 ss.n341 ss.n340 8.75769
R386 ss.n117 ss.n116 8.63854
R387 ss.n199 ss.n198 8.6074
R388 ss.n313 ss.n312 8.40926
R389 ss.n172 ring_100mV_0.SS 8.05129
R390 ss.n291 ss.t40 6.97557
R391 ss.n178 ss.n177 6.963
R392 ss.n0 ss.t67 6.96143
R393 ss.n1 ss.t66 6.96143
R394 ss.n198 ss.t85 6.96143
R395 ss.n196 ss.t84 6.96143
R396 ss.n13 ss.t90 6.96143
R397 ss.n4 ss.t91 6.96143
R398 ss.n186 ss.t81 6.96143
R399 ss.n48 ss.t80 6.96143
R400 ss.n238 ss.n226 6.73922
R401 ss.n134 ss.n131 6.32011
R402 ss.n368 ss.n367 5.9778
R403 ss.n373 ss.n372 5.9778
R404 ss.n59 ss.t167 5.95384
R405 ss.n52 ss.t132 5.95384
R406 ss.n152 ss.t129 5.86529
R407 ss.n149 ss.t163 5.86456
R408 iref_2nA_0.iref_2nA_mirrors_0.SS ss.n439 5.6745
R409 ss.n326 ss.n325 5.36738
R410 ss.n327 ss.n326 5.36738
R411 ss.n328 ss.n327 5.21979
R412 ss.n314 ss.n311 5.2134
R413 ring_100mV_0.mdls_inv_3.SS ss.n148 5.21317
R414 ss.n314 ss.n313 5.16179
R415 ss.n83 ring_100mV_0.mdls_inv_5.SS 5.1001
R416 ss.n267 ring_100mV_0.mdls_inv_7.SS 5.1001
R417 ss.n360 ring_100mV_0.mdls_inv_9.SS 5.1001
R418 ss.n345 ring_100mV_0.mdls_inv_0.SS 5.1001
R419 ss.n141 ss.n69 5.04939
R420 ss.n337 ldo_0.SS 4.99932
R421 ss.n441 ss.n440 4.93732
R422 ss.n163 ss.n162 4.80538
R423 ss.n72 ss.n71 4.80538
R424 ss.n59 ss.t226 4.59778
R425 ss.n60 ss.t217 4.59778
R426 ss.n52 ss.t7 4.59778
R427 ss.n53 ss.t198 4.59778
R428 ss.n54 ss.t224 4.59778
R429 ss.n61 ss.t211 4.55016
R430 ss.n62 ss.t114 4.55016
R431 ss.n63 ss.t53 4.55016
R432 ss.n64 ss.t118 4.55016
R433 ss.n65 ss.t231 4.55016
R434 ss.n58 ss.t104 4.55016
R435 ss.n57 ss.t229 4.55016
R436 ss.n56 ss.t46 4.55016
R437 ss.n55 ss.t100 4.55016
R438 ss.n152 ss.t22 4.50985
R439 ss.n149 ss.t108 4.5085
R440 ss.n150 ss.t39 4.46515
R441 ss.n151 ss.t137 4.4579
R442 ss.n154 ss.t5 4.4579
R443 ss.n153 ss.t173 4.4579
R444 ss.n352 ss.n292 4.43918
R445 ss.n16 ss.n13 4.35124
R446 ss.n206 ss 4.30941
R447 ss.n430 ss 4.2532
R448 ring_100mV_0.SS ss.n170 4.14018
R449 ss.n87 ss.n85 4.09668
R450 ss.n264 ss.n263 4.09668
R451 ss.n363 ss.n362 4.09668
R452 ss.n342 ss.n341 4.09668
R453 ss.n331 ss.n257 4.09668
R454 ss.n384 ss.n383 4.09668
R455 ss.n397 ss.n396 4.09668
R456 ss.n419 ss.n418 4.09668
R457 ss.n248 ss.n247 4.09668
R458 ss.n256 ss.n255 4.09668
R459 ss.t177 ss.t9 3.98691
R460 ss.t192 ss.t171 3.98691
R461 ss.t44 ss.t130 3.98691
R462 ss.t232 ss.t127 3.98691
R463 ss.t98 ss.t161 3.98691
R464 ss.t181 ss.t13 3.89258
R465 ss.t206 ss.t10 3.89258
R466 ss.t30 ss.t200 3.89258
R467 ss.t35 ss.t151 3.89258
R468 ss.t155 ss.t146 3.89258
R469 ss.n319 ss.t74 3.41269
R470 ss.n329 ss.t95 3.41269
R471 ss.n373 ss.t196 3.16453
R472 ss.n246 ss.t111 3.16453
R473 ss.n408 ss.t194 3.16453
R474 ss.n399 ss.t43 3.16453
R475 ss.n382 ss.t189 3.16453
R476 ss.n83 ss.t186 3.16453
R477 ss.n267 ss.t19 3.16453
R478 ss.n360 ss.t202 3.16453
R479 ss.n345 ss.t27 3.16453
R480 ss.n367 ss.t150 3.16453
R481 ss.n170 ring_100mV_0.SS 3.14741
R482 ss.n322 ss.n321 3.09416
R483 ss.n436 ss.n203 2.99115
R484 ss.n388 ss.n378 2.99081
R485 ss.n406 ss.n402 2.99081
R486 ss.n414 ss.n411 2.99081
R487 ss.n252 ss.n242 2.99081
R488 ss.n80 ss.n79 2.92006
R489 ss.n272 ss.n262 2.92006
R490 ss.n357 ss.n356 2.92006
R491 ss.n350 ss.n293 2.92006
R492 ss.n325 ss.n324 2.8852
R493 ss.n440 iref_2nA_0.iref_2nA_mirrors_0.SS 2.81516
R494 ss.n194 ss.n192 2.69854
R495 iref_2nA_0.SS ss.n47 2.52476
R496 iref_2nA_0.SS ss.n441 2.48008
R497 ss.n429 ss.n424 2.3819
R498 ss.n116 ss.n115 2.2502
R499 ss.n169 ss.n161 2.24002
R500 ss.n183 ss.n178 2.20466
R501 ldo_0.SS ss.n336 1.74251
R502 ss.n188 ss.n187 1.601
R503 ss.n334 ss.n329 1.38918
R504 ss.n150 ss.n149 1.37246
R505 ss.n60 ss.n59 1.35656
R506 ss.n53 ss.n52 1.35656
R507 ss.n54 ss.n53 1.35656
R508 ss.n61 ss.n60 1.33075
R509 ss.n189 ss.n188 1.28727
R510 ss.n36 ss.n35 1.24652
R511 ss.n95 ss.n94 1.13695
R512 ss.n230 ss.n229 1.08301
R513 ss.n203 ss.n199 0.997385
R514 ss.n320 ss.n319 0.989591
R515 ss.t93 ss.t152 0.973521
R516 ss.n232 ss.n227 0.945812
R517 ss.n235 ss.n234 0.945812
R518 ss.n55 ss.n54 0.915706
R519 ss.n161 ss.n158 0.753441
R520 ss.n236 ss.n235 0.594703
R521 ss.n232 ss.n231 0.585645
R522 ss.n233 ss.n232 0.58021
R523 ss.n235 ss.n233 0.571152
R524 ss.n226 ss.n215 0.57063
R525 ss.n93 ss.n90 0.569131
R526 ss.n137 ss.n136 0.500622
R527 ss.n237 ss.n236 0.441037
R528 ss.n323 ss.n322 0.387207
R529 ss.n154 ss.n153 0.329447
R530 ss.n151 ss.n150 0.329292
R531 ss.n153 ss.n152 0.316559
R532 ss.n155 ss.n151 0.307243
R533 ss.n319 ss.n318 0.291409
R534 ss.n231 ss.n230 0.254123
R535 ss.n56 ss.n55 0.238595
R536 ss.n57 ss.n56 0.238595
R537 ss.n58 ss.n57 0.238595
R538 ss.n65 ss.n64 0.238595
R539 ss.n64 ss.n63 0.238595
R540 ss.n63 ss.n62 0.238595
R541 ss.n62 ss.n61 0.238595
R542 ss.n226 ss.n225 0.190812
R543 ss.n66 ss.n58 0.18919
R544 ss.n238 ss.n237 0.139656
R545 ss.n229 ss.n228 0.0932419
R546 ss.n172 ss.n171 0.0766905
R547 ss.n135 ss.n134 0.0499686
R548 ss.n66 ss.n65 0.0499048
R549 ss.n23 ss.n22 0.0425017
R550 ss.n22 ss.n21 0.0425017
R551 ss.n206 ss.n205 0.0425017
R552 ss.n205 ss.n204 0.0425017
R553 ss.n287 ss.n286 0.0360926
R554 ss.n288 ss.n287 0.0360926
R555 ss.n339 ss.n338 0.0360926
R556 ss.n340 ss.n339 0.0360926
R557 ss.n155 ss.n154 0.0227039
R558 ss.n27 ss.n26 0.0128626
R559 ss.t62 ss.n27 0.0128626
R560 ss.t62 ss.n19 0.0128626
R561 ss.n19 ss.n18 0.0128626
R562 ss.n290 ss.n289 0.00609809
R563 ss.n291 ss.n290 0.00609809
R564 ss.n284 ss.n283 0.00609809
R565 ss.n283 ss.n282 0.00609809
R566 ss.n121 ss.n120 0.00358142
R567 ss.n122 ss.n121 0.00233142
R568 ss.n356 ss.n354 0.00200294
R569 ss.n272 ss.n270 0.00200294
R570 ss.n79 ss.n76 0.00200294
R571 ss.n350 ss.n348 0.00200294
R572 ss.n387 ss.n386 0.00200294
R573 ss.n405 ss.n404 0.00200294
R574 ss.n416 ss.n415 0.00200294
R575 ss.n251 ss.n250 0.00200294
R576 ss.n93 ss.n92 0.00150773
R577 ss.n94 ss.n93 0.00150002
R578 ss.n215 ss.n214 0.00107233
R579 ss.n120 ss.n118 0.00101107
R580 ss.n120 ss.n119 0.0010106
R581 ss.n343 ss.n293 0.00100729
R582 ss.n358 ss.n357 0.00100729
R583 ss.n265 ss.n262 0.00100729
R584 ss.n81 ss.n80 0.00100729
R585 ss.n92 ss.n91 0.00100729
R586 ss.n380 ss.n378 0.00100728
R587 ss.n402 ss.n401 0.00100728
R588 ss.n411 ss.n410 0.00100728
R589 ss.n244 ss.n242 0.00100728
R590 ss.n160 ss.n159 0.00100728
R591 ss.n344 ss.n343 0.00100728
R592 ss.n359 ss.n358 0.00100728
R593 ss.n266 ss.n265 0.00100728
R594 ss.n82 ss.n81 0.00100728
R595 ss.n381 ss.n380 0.00100728
R596 ss.n401 ss.n400 0.00100728
R597 ss.n410 ss.n409 0.00100728
R598 ss.n245 ss.n244 0.00100728
R599 ss.n224 ss.n221 0.00100463
R600 ss.n76 ss.n75 0.00100294
R601 ss.n270 ss.n269 0.00100294
R602 ss.n354 ss.n353 0.00100294
R603 ss.n388 ss.n387 0.00100294
R604 ss.n406 ss.n405 0.00100294
R605 ss.n415 ss.n414 0.00100294
R606 ss.n252 ss.n251 0.00100294
R607 ss.n348 ss.n347 0.00100294
R608 ss.n217 ss.n216 0.000530441
R609 ss.n10 ss.n9 0.000524964
R610 ss.n9 ss.n8 0.000524964
R611 ss.n174 ss.n173 0.000524415
R612 ss.n175 ss.n174 0.000524415
R613 ss.n177 ss.n176 0.000519599
R614 ss.n212 ss.n211 0.000518216
R615 ss.n211 ss.n210 0.000518216
R616 ss.n203 ss.n202 0.000518064
R617 ss.n202 ss.n201 0.000518064
R618 ss.n16 ss.n15 0.000518064
R619 ss.n15 ss.n14 0.000518064
R620 ss.n440 ss.n51 0.000518064
R621 ss.n51 ss.n50 0.000518064
R622 ss.n34 ss.n33 0.000518064
R623 ss.n33 ss.n32 0.000518064
R624 ss.n350 ss.n349 0.000513494
R625 ss.n356 ss.n355 0.000513494
R626 ss.n272 ss.n271 0.000513494
R627 ss.n79 ss.n78 0.000513494
R628 ss.n90 ss.n89 0.000513494
R629 ss.n169 ss.n168 0.000513494
R630 ss.n168 ss.n167 0.000513494
R631 ss.n388 ss.n379 0.000513494
R632 ss.n406 ss.n403 0.000513494
R633 ss.n414 ss.n413 0.000513494
R634 ss.n252 ss.n243 0.000513494
R635 ss.n140 ss.n139 0.000513051
R636 ss.n139 ss.n138 0.000513051
R637 ss.n318 ss.n317 0.00051152
R638 ss.n317 ss.n316 0.00051152
R639 ss.n334 ss.n333 0.00051152
R640 ss.n333 ss.n332 0.00051152
R641 ss.n46 ss.n45 0.000511457
R642 ss.n45 ss.n44 0.000511457
R643 ss.n118 ss.n117 0.00051107
R644 ss.n131 ss.n130 0.000510324
R645 ss.n130 ss.n129 0.000510324
R646 ss.n280 ss.n279 0.000510263
R647 ss.n279 ss.n278 0.000510263
R648 ss.n110 ss.n109 0.000510194
R649 ss.n126 ss.n110 0.000510194
R650 ss.n125 ss.n124 0.000510194
R651 ss.n126 ss.n125 0.000510194
R652 ss.n161 ss.n160 0.00050775
R653 ss.n30 ss.n29 0.000506779
R654 ss.n29 ss.n28 0.000506779
R655 ss.n42 ss.n41 0.000505267
R656 ss.n43 ss.n42 0.000505267
R657 ss.n221 ss.n220 0.000504934
R658 ss.n241 ss.n240 0.000504379
R659 ss.n240 ss.n239 0.000504379
R660 ss.n100 ss.n99 0.000504346
R661 ss.n99 ss.n98 0.000504346
R662 ss.n300 ss.n299 0.000503106
R663 ss.n301 ss.n300 0.000503106
R664 ss.n303 ss.n302 0.000503106
R665 ss.n302 ss.n301 0.000503106
R666 ss.n74 ss.n73 0.000502943
R667 ss.n89 ss.n74 0.000502943
R668 ss.n165 ss.n164 0.000502943
R669 ss.n167 ss.n165 0.000502943
R670 ss.n277 ss.n276 0.000502681
R671 ss.n276 ss.n275 0.000502681
R672 ss.n147 ss.n146 0.000502057
R673 ss.n146 ss.n145 0.000502057
R674 ss.n310 ss.n309 0.000501887
R675 ss.n309 ss.n308 0.000501887
R676 ss.n105 ss.n104 0.00050184
R677 ss.n104 ss.n103 0.00050184
R678 ss.n182 ss.n181 0.00050184
R679 ss.n181 ss.n180 0.00050184
R680 ss.n142 ss.n141 0.000501833
R681 ss.n143 ss.n142 0.000501833
R682 ss.n371 ss.n370 0.000501787
R683 ss.n370 ss.n369 0.000501787
R684 ss.n128 ss.n127 0.000501613
R685 ss.n127 ss.n126 0.000501613
R686 ss.n108 ss.n107 0.000501613
R687 ss.n107 ss.n106 0.000501613
R688 ss.n134 ss.n133 0.000501511
R689 ss.n133 ss.n132 0.000501511
R690 ss.n115 ss.n114 0.000501511
R691 ss.n114 ss.n113 0.000501511
R692 ss.n429 ss.n428 0.000501075
R693 ss.n428 ss.n427 0.000501075
R694 ss.n392 ss.n391 0.000501075
R695 ss.n391 ss.n390 0.000501075
R696 ss.n365 ss.n364 0.000500622
R697 ss.n422 ss.n421 0.000500622
R698 ss.n421 ss.n420 0.000500622
R699 ss.n435 ss.n434 0.000500587
R700 ss.n434 ss.n433 0.000500587
R701 ss.n394 ss.n393 0.000500387
R702 ss.n395 ss.n394 0.000500387
R703 ss.n158 ss.n157 0.000500208
R704 ss.n157 ss.n156 0.000500208
R705 ss.n69 ss.n68 0.000500141
R706 ss.n68 ss.n67 0.000500141
R707 ss.n158 ss.n155 0.000500116
R708 ss.n69 ss.n66 0.000500044
R709 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t22 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t19 75.728
R710 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t13 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t22 75.728
R711 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t17 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t13 75.728
R712 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t24 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t17 75.728
R713 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t12 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t24 75.728
R714 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t14 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t12 75.728
R715 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t20 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t14 75.728
R716 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t25 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t20 75.728
R717 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t16 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t25 75.728
R718 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t21 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t16 75.728
R719 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t23 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t21 75.728
R720 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t15 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t23 75.728
R721 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n6 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t18 37.8646
R722 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n6 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t15 37.8639
R723 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n4 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t11 12.8247
R724 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n5 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t8 12.8247
R725 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n2 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t7 12.8247
R726 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n3 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t3 12.8247
R727 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n0 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t6 11.428
R728 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n4 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t1 11.428
R729 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n5 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t2 11.428
R730 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n1 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t9 11.428
R731 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n2 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t10 11.428
R732 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n3 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t0 11.428
R733 iref_2nA_0.iref_2nA_mirrors_0.Ip2 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n1 8.50055
R734 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n7 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t5 8.17164
R735 iref_2nA_0.iref_2nA_igenerator_0.Ip2 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t4 7.50959
R736 iref_2nA_0.iref_2nA_mirrors_0.Ip2 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n7 5.32175
R737 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n7 iref_2nA_0.iref_2nA_igenerator_0.Ip2 3.49672
R738 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n0 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n6 2.74398
R739 iref_2nA_0.iref_2nA_mirrors_0.Ip2 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n0 0.990509
R740 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n0 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n5 0.810482
R741 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n1 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n3 0.810433
R742 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n0 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n4 0.810432
R743 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n1 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n2 0.810432
R744 a_1555_7968.n0 a_1555_7968.t3 37.8394
R745 a_1555_7968.n0 a_1555_7968.t1 37.8394
R746 a_1555_7968.t0 a_1555_7968.n0 12.0988
R747 a_1555_7968.n0 a_1555_7968.t2 11.4337
R748 a_1555_7968.n0 a_1555_7968.t5 11.428
R749 a_1555_7968.n0 a_1555_7968.t4 11.428
R750 dd_01.n26 dd_01.n25 7521.18
R751 dd_01.n32 dd_01.n26 7517.65
R752 dd_01.n30 dd_01.n25 7517.65
R753 dd_01.n32 dd_01.n30 7514.12
R754 dd_01.n21 dd_01.n20 2985.88
R755 dd_01.n18 dd_01.n16 2985.88
R756 dd_01.n16 dd_01.n15 949.587
R757 dd_01.n20 dd_01.n19 949.587
R758 dd_01.n139 dd_01.n134 622.683
R759 dd_01.n29 dd_01.n27 459.671
R760 dd_01.n29 dd_01.n28 452.519
R761 dd_01.n137 dd_01.t2 431.565
R762 dd_01.t74 dd_01.t55 367.363
R763 dd_01.t26 dd_01.t74 367.363
R764 dd_01.t29 dd_01.t35 367.363
R765 dd_01.t65 dd_01.t29 367.363
R766 dd_01.n149 dd_01.n148 344.031
R767 dd_01.n137 dd_01.t33 319.678
R768 dd_01.n17 dd_01.n13 318.495
R769 dd_01.n17 dd_01.n14 318.495
R770 dd_01.n22 dd_01.n14 282.247
R771 dd_01.n11 dd_01.n8 243.716
R772 dd_01.t55 dd_01.n25 232.912
R773 dd_01.n143 dd_01.n132 226.184
R774 dd_01.n32 dd_01.t65 213.075
R775 dd_01.n23 dd_01.n13 209.695
R776 dd_01.n11 dd_01.n10 208.559
R777 dd_01.t1 dd_01.n127 202.427
R778 dd_01.n47 dd_01.t18 199.849
R779 dd_01.t35 dd_01.n31 193.233
R780 dd_01.n146 dd_01.t1 192.995
R781 dd_01.n143 dd_01.n139 189.365
R782 dd_01.n31 dd_01.t26 174.131
R783 dd_01.n5 dd_01.n2 157.536
R784 dd_01.t24 dd_01.n73 119.335
R785 dd_01.n89 dd_01.t22 96.026
R786 dd_01.n101 dd_01.t44 89.4352
R787 dd_01.n103 dd_01.t43 89.4352
R788 dd_01.n120 dd_01.t59 89.4352
R789 dd_01.n55 dd_01.t50 89.4352
R790 dd_01.n62 dd_01.t63 89.4352
R791 dd_01.n33 dd_01.n27 89.3686
R792 dd_01.n89 dd_01.t24 67.1251
R793 dd_01.n92 dd_01.n65 62.6718
R794 dd_01.n92 dd_01.n63 62.6718
R795 dd_01.n27 dd_01.t67 60.0995
R796 dd_01.n28 dd_01.t57 60.0995
R797 dd_01.t0 dd_01.n116 59.4732
R798 dd_01.n52 dd_01.n51 58.4844
R799 dd_01.n51 dd_01.n50 58.4844
R800 dd_01.n110 dd_01.n109 58.4844
R801 dd_01.n111 dd_01.n110 58.4844
R802 dd_01.n112 dd_01.n111 58.4844
R803 dd_01.n108 dd_01.n107 58.4844
R804 dd_01.n107 dd_01.n106 58.4844
R805 dd_01.n57 dd_01.n56 58.4844
R806 dd_01.n58 dd_01.n57 58.4844
R807 dd_01.n59 dd_01.n58 58.4844
R808 dd_01.t3 dd_01.n114 58.3834
R809 dd_01.n122 dd_01.t60 57.7693
R810 dd_01.n60 dd_01.t62 57.1406
R811 dd_01.n53 dd_01.t49 57.1406
R812 dd_01.n74 dd_01.t73 57.1406
R813 dd_01.n75 dd_01.t72 57.1406
R814 dd_01.n82 dd_01.t47 57.1406
R815 dd_01.n81 dd_01.t46 57.1406
R816 dd_01.n66 dd_01.t52 57.1406
R817 dd_01.n67 dd_01.t53 57.1406
R818 dd_01.n63 dd_01.t40 57.1406
R819 dd_01.n65 dd_01.t41 57.1406
R820 dd_01.n128 dd_01.t70 57.1406
R821 dd_01.n54 dd_01.n53 53.2677
R822 dd_01.n34 dd_01.n33 49.5403
R823 dd_01.n122 dd_01.n121 44.9447
R824 dd_01.n53 dd_01.n52 44.2622
R825 dd_01.n60 dd_01.n59 44.2622
R826 dd_01.n24 dd_01.n23 41.6985
R827 dd_01.n92 dd_01.n91 41.2005
R828 dd_01.n131 dd_01.n129 40.1187
R829 dd_01.n124 dd_01.n122 39.5995
R830 dd_01.n94 dd_01.n93 38.9913
R831 dd_01.n100 dd_01.n99 38.8928
R832 dd_01.n99 dd_01.n98 38.8928
R833 dd_01.n100 dd_01.n92 38.282
R834 dd_01.n40 dd_01.n39 34.174
R835 dd_01.n39 dd_01.n38 34.174
R836 dd_01.n36 dd_01.n35 34.174
R837 dd_01.n35 dd_01.n34 34.174
R838 dd_01.n34 dd_01.t66 32.0995
R839 dd_01.n35 dd_01.t30 32.0995
R840 dd_01.n36 dd_01.t36 32.0995
R841 dd_01.n38 dd_01.t27 32.0995
R842 dd_01.n39 dd_01.t75 32.0995
R843 dd_01.n40 dd_01.t56 32.0995
R844 dd_01.n113 dd_01.n112 30.1336
R845 dd_01.n113 dd_01.n108 28.3513
R846 dd_01.n117 dd_01.t3 28.2824
R847 dd_01.n117 dd_01.t0 27.6433
R848 dd_01.n77 dd_01.n75 26.9918
R849 dd_01.n80 dd_01.n74 26.9918
R850 dd_01.n86 dd_01.n81 26.9918
R851 dd_01.n83 dd_01.n82 26.9918
R852 dd_01.n68 dd_01.n67 26.9918
R853 dd_01.n71 dd_01.n66 26.9918
R854 dd_01.n41 dd_01.n40 26.4458
R855 dd_01.n93 dd_01.t32 25.9683
R856 dd_01.n94 dd_01.t23 25.9683
R857 dd_01.n98 dd_01.t25 25.9683
R858 dd_01.n99 dd_01.t31 25.9683
R859 dd_01.n61 dd_01.n60 25.6869
R860 dd_01.t33 dd_01.t69 25.0188
R861 dd_01.n121 dd_01.n120 22.1276
R862 dd_01.n55 dd_01.n54 22.1276
R863 dd_01.n87 dd_01.n80 22.124
R864 iref_2nA_0.iref_2nA_vref_0.DD dd_01.n142 22.0801
R865 dd_01.n125 dd_01.n124 21.3338
R866 dd_01.n97 dd_01.n94 19.5943
R867 dd_01.n98 dd_01.n97 19.0036
R868 dd_01.n37 dd_01.n36 18.0327
R869 dd_01.n77 dd_01.n76 17.0289
R870 dd_01.n132 dd_01.n131 16.7789
R871 dd_01.n38 dd_01.n37 16.1418
R872 dd_01.n119 dd_01.n55 16.1067
R873 dd_01.n103 dd_01.n102 15.5135
R874 dd_01.n102 dd_01.n101 15.5135
R875 dd_01.n62 dd_01.n61 15.5135
R876 dd_01.n120 dd_01.n119 15.0827
R877 dd_01.n79 dd_01.n77 14.4898
R878 dd_01.n80 dd_01.n79 14.4898
R879 dd_01.n86 dd_01.n85 14.4898
R880 dd_01.n85 dd_01.n83 14.4898
R881 dd_01.n102 dd_01.t42 13.7387
R882 dd_01.n61 dd_01.t61 13.7387
R883 dd_01.n54 dd_01.t48 13.7387
R884 dd_01.n121 dd_01.t58 13.7387
R885 dd_01.n79 dd_01.t71 13.7387
R886 dd_01.t71 dd_01.n78 13.7387
R887 dd_01.n85 dd_01.t45 13.7387
R888 dd_01.t45 dd_01.n84 13.7387
R889 dd_01.n70 dd_01.t51 13.7387
R890 dd_01.t51 dd_01.n69 13.7387
R891 dd_01.n92 dd_01.t39 13.7387
R892 dd_01.t39 dd_01.n64 13.7387
R893 dd_01.n71 dd_01.n70 13.7236
R894 dd_01.n70 dd_01.n68 13.7236
R895 dd_01.n125 dd_01.n49 13.177
R896 dd_01.n132 dd_01.t34 12.0543
R897 dd_01.n45 dd_01.t20 11.8558
R898 dd_01.n49 dd_01.t19 11.4275
R899 dd_01.n59 dd_01.t10 11.4275
R900 dd_01.n58 dd_01.t7 11.4275
R901 dd_01.n57 dd_01.t16 11.4275
R902 dd_01.n56 dd_01.t12 11.4275
R903 dd_01.n106 dd_01.t5 11.4275
R904 dd_01.n107 dd_01.t17 11.4275
R905 dd_01.n108 dd_01.t15 11.4275
R906 dd_01.n112 dd_01.t9 11.4275
R907 dd_01.n111 dd_01.t4 11.4275
R908 dd_01.n110 dd_01.t13 11.4275
R909 dd_01.n109 dd_01.t8 11.4275
R910 dd_01.n50 dd_01.t6 11.4275
R911 dd_01.n51 dd_01.t14 11.4275
R912 dd_01.n52 dd_01.t11 11.4275
R913 dd_01.n101 dd_01.n100 10.6672
R914 iref_2nA_0.DD dd_01.n154 10.2882
R915 dd_01.n104 dd_01.n62 9.82907
R916 dd_01.n41 dd_01.t54 9.47999
R917 dd_01.n33 dd_01.t64 9.47999
R918 dd_01.n104 dd_01.n103 9.21955
R919 dd_01.n154 dd_01.n46 8.85536
R920 dd_01.n143 iref_2nA_0.iref_2nA_vref_0.DD 8.72328
R921 dd_01.n42 dd_01.n24 7.69412
R922 dd_01.n87 dd_01.n86 6.71433
R923 dd_01.n28 dd_01.n24 6.51432
R924 dd_01.n91 dd_01.n71 5.61588
R925 dd_01.n22 dd_01.t38 5.52608
R926 dd_01.n42 dd_01.n41 5.23543
R927 dd_01.n0 dd_01.t28 4.89002
R928 dd_01.n0 dd_01.t21 4.38996
R929 dd_01.n154 dd_01.n153 4.28102
R930 dd_01.n43 dd_01.n12 4.17205
R931 dd_01.n128 dd_01.t68 4.11799
R932 dd_01.n154 dd_01.n45 3.99011
R933 dd_01.n153 dd_01 2.82647
R934 iref_2nA_0.DD dd_01.n44 2.56417
R935 dd_01.n144 dd_01.n143 2.44683
R936 dd_01.n44 dd_01.n43 2.42546
R937 dd_01.n23 dd_01.n22 1.98969
R938 dd_01.n129 dd_01.n128 1.54124
R939 ldo_0.DD dd_01.n42 1.39885
R940 dd_01.n149 dd_01.n125 0.970197
R941 dd_01.n44 dd_01 0.861062
R942 dd_01.n124 dd_01.n123 0.706994
R943 dd_01.n123 dd_01 0.644656
R944 dd_01.n43 ldo_0.DD 0.464881
R945 dd_01.n142 dd_01.n141 0.332968
R946 dd_01.n48 dd_01.n47 0.28389
R947 dd_01.n12 vref01_0.DD 0.0698807
R948 dd_01.n141 dd_01.n140 0.0402849
R949 dd_01.n140 dd_01.n48 0.0402849
R950 dd_01.n16 dd_01.n13 0.025954
R951 dd_01.n20 dd_01.n14 0.025954
R952 vref01_0.DD dd_01.n0 0.0182752
R953 dd_01.n151 dd_01.n150 0.0146429
R954 dd_01.n150 dd_01.n149 0.0141431
R955 dd_01.n5 dd_01.n4 0.00768538
R956 dd_01.n7 dd_01.n6 0.0076851
R957 dd_01.n8 dd_01.n7 0.00740969
R958 dd_01.n4 dd_01.n3 0.00740969
R959 dd_01.n152 dd_01.n151 0.00674884
R960 dd_01.n153 dd_01.n152 0.00624891
R961 dd_01.n33 dd_01.n32 0.00450849
R962 dd_01.n41 dd_01.n25 0.00450849
R963 dd_01.n134 dd_01.n133 0.00424858
R964 dd_01.n131 dd_01.n130 0.00424858
R965 dd_01.n18 dd_01.n17 0.00414317
R966 dd_01.n22 dd_01.n21 0.00414317
R967 dd_01.n145 dd_01.n144 0.00377503
R968 dd_01.n146 dd_01.n145 0.00377503
R969 dd_01.n147 dd_01.n146 0.00377503
R970 dd_01.n148 dd_01.n147 0.00377503
R971 dd_01.n119 dd_01.n118 0.00369903
R972 dd_01.n118 dd_01.n117 0.00369903
R973 dd_01.n105 dd_01.n104 0.00369903
R974 dd_01.n117 dd_01.n105 0.00369903
R975 dd_01.n21 dd_01.n15 0.00355895
R976 dd_01.n19 dd_01.n18 0.00348454
R977 dd_01.n88 dd_01.n87 0.00338999
R978 dd_01.n89 dd_01.n88 0.00338999
R979 dd_01.n90 dd_01.n89 0.00338999
R980 dd_01.n91 dd_01.n90 0.00338999
R981 dd_01.n127 dd_01.n126 0.00337446
R982 dd_01.n2 dd_01.n1 0.00271961
R983 dd_01.n10 dd_01.n9 0.00271961
R984 dd_01.n136 dd_01.n135 0.00268001
R985 dd_01.n137 dd_01.n136 0.00268001
R986 dd_01.n139 dd_01.n138 0.00268001
R987 dd_01.n138 dd_01.n137 0.00268001
R988 dd_01.t37 dd_01.n15 0.00231816
R989 dd_01.n19 dd_01.t37 0.00215862
R990 dd_01.n37 dd_01.n26 0.00193193
R991 dd_01.n31 dd_01.n26 0.00193193
R992 dd_01.n31 dd_01.n30 0.00193193
R993 dd_01.n30 dd_01.n29 0.00193193
R994 dd_01.n73 dd_01.n72 0.00161095
R995 dd_01.n97 dd_01.n96 0.00161095
R996 dd_01.n96 dd_01.n95 0.00161095
R997 dd_01.n6 dd_01.t76 0.00122457
R998 dd_01.t76 dd_01.n5 0.0012243
R999 dd_01.n151 dd_01.n48 0.00100005
R1000 dd_01.n12 dd_01.n11 0.00094942
R1001 dd_01.n114 dd_01.n113 0.000866167
R1002 dd_01.n116 dd_01.n115 0.000866167
R1003 dd_02.n162 dd_02.n157 4743.53
R1004 dd_02.n177 dd_02.n157 4740
R1005 dd_02.n162 dd_02.n158 4740
R1006 dd_02.n177 dd_02.n158 4736.47
R1007 dd_02.n174 dd_02.n164 3331.76
R1008 dd_02.n174 dd_02.n165 3331.76
R1009 dd_02.n170 dd_02.n164 3331.76
R1010 dd_02.n170 dd_02.n165 3331.76
R1011 dd_02.n161 dd_02.n159 505.976
R1012 dd_02.n159 dd_02.n156 487.529
R1013 dd_02.n161 dd_02.n160 450.673
R1014 dd_02.t20 dd_02.t16 380.762
R1015 dd_02.t24 dd_02.t22 380.762
R1016 dd_02.n171 dd_02.n168 355.389
R1017 dd_02.n168 dd_02.n166 354.635
R1018 dd_02.n175 dd_02.t41 353.156
R1019 dd_02.n170 dd_02.t0 351.26
R1020 dd_02.n173 dd_02.n172 345.601
R1021 dd_02.n172 dd_02.n171 345.601
R1022 dd_02.n176 dd_02.t24 318.889
R1023 dd_02.t16 dd_02.n162 317.942
R1024 dd_02.n85 dd_02.t40 223.291
R1025 dd_02.n41 dd_02.t37 223.291
R1026 dd_02.n54 dd_02.t10 223.291
R1027 dd_02.n29 dd_02.t31 223.291
R1028 dd_02.n6 dd_02.t18 223.291
R1029 dd_02.n31 dd_02.t32 223.291
R1030 dd_02.n60 dd_02.t11 223.291
R1031 dd_02.n47 dd_02.t34 223.291
R1032 dd_02.n70 dd_02.t27 223.291
R1033 dd_02.n19 dd_02.t7 223.291
R1034 dd_02.n179 dd_02.n178 192.433
R1035 dd_02.n163 dd_02.t20 191.333
R1036 dd_02.t0 dd_02.n169 191.333
R1037 dd_02.t22 dd_02.n163 189.429
R1038 dd_02.n169 dd_02.t41 189.429
R1039 dd_02.n43 dd_02.n42 156.236
R1040 dd_02.n56 dd_02.n55 156.236
R1041 dd_02.n99 dd_02.n30 156.236
R1042 dd_02.n135 dd_02.n7 156.236
R1043 dd_02.n95 dd_02.n32 156.236
R1044 dd_02.n62 dd_02.n61 156.236
R1045 dd_02.n49 dd_02.n48 156.236
R1046 dd_02.n72 dd_02.n71 156.236
R1047 dd_02.n21 dd_02.n20 152.847
R1048 dd_02.n87 dd_02.n86 151.719
R1049 dd_02.n179 dd_02.n155 150.099
R1050 dd_02.n176 dd_02.n175 145.642
R1051 dd_02.n85 dd_02.t3 133.543
R1052 dd_02.n41 dd_02.t39 133.543
R1053 dd_02.n54 dd_02.t9 133.543
R1054 dd_02.n29 dd_02.t29 133.543
R1055 dd_02.n6 dd_02.t28 133.543
R1056 dd_02.n31 dd_02.t26 133.543
R1057 dd_02.n60 dd_02.t12 133.543
R1058 dd_02.n47 dd_02.t36 133.543
R1059 dd_02.n70 dd_02.t19 133.543
R1060 dd_02.n19 dd_02.t4 133.543
R1061 dd_02.n172 dd_02.n167 78.0313
R1062 ring_100mV_0.mdls_inv_5.DD dd_02.n43 72.0212
R1063 ring_100mV_0.mdls_inv_7.DD dd_02.n56 72.0212
R1064 dd_02.n99 ring_100mV_0.mdls_inv_9.DD 72.0212
R1065 dd_02 dd_02.n135 72.0212
R1066 ring_100mV_0.mdls_inv_8.DD dd_02.n95 67.8992
R1067 dd_02.n62 ring_100mV_0.mdls_inv_6.DD 67.8992
R1068 dd_02.n49 ring_100mV_0.mdls_inv_4.DD 67.8992
R1069 dd_02.n72 ring_100mV_0.mdls_inv_1.DD 67.8992
R1070 dd_02.n138 dd_02.n137 66.1197
R1071 dd_02.n97 dd_02.n96 66.1197
R1072 dd_02.n58 dd_02.n57 66.1197
R1073 dd_02.n45 dd_02.n44 66.1197
R1074 dd_02.n36 ring_100mV_0.mdls_inv_3.DD 65.5729
R1075 dd_02.n167 dd_02.t1 65.041
R1076 dd_02.n143 dd_02.n142 64.9329
R1077 dd_02.n167 dd_02.t42 64.529
R1078 dd_02.n138 dd_02.n136 62.5594
R1079 dd_02.n98 dd_02.n97 62.5594
R1080 dd_02.n59 dd_02.n58 62.5594
R1081 dd_02.n46 dd_02.n45 62.5594
R1082 dd_02.n86 dd_02.n85 60.6614
R1083 dd_02.n42 dd_02.n41 60.6614
R1084 dd_02.n55 dd_02.n54 60.6614
R1085 dd_02.n30 dd_02.n29 60.6614
R1086 dd_02.n7 dd_02.n6 60.6614
R1087 dd_02.n32 dd_02.n31 60.6614
R1088 dd_02.n61 dd_02.n60 60.6614
R1089 dd_02.n48 dd_02.n47 60.6614
R1090 dd_02.n71 dd_02.n70 60.6614
R1091 dd_02.n20 dd_02.n19 60.6614
R1092 dd_02.n23 dd_02.n18 31.5911
R1093 dd_02.n89 dd_02.n84 31.249
R1094 dd_02.n153 dd_02.t17 30.1358
R1095 dd_02.n154 dd_02.t25 30.1029
R1096 dd_02.n152 dd_02.t21 28.8743
R1097 dd_02.n152 dd_02.t23 28.8743
R1098 dd_02.n24 dd_02.t35 28.5685
R1099 dd_02.n38 dd_02.t33 28.5685
R1100 dd_02.n128 dd_02.t6 28.5685
R1101 dd_02.n125 dd_02.t38 28.5685
R1102 dd_02.n122 dd_02.t8 28.5685
R1103 dd_02.n119 dd_02.t30 28.5685
R1104 dd_02.n67 dd_02.t15 28.5685
R1105 dd_02.n64 dd_02.t13 28.5685
R1106 dd_02.n51 dd_02.t14 28.5685
R1107 dd_02.n90 dd_02.t43 28.5685
R1108 dd_02.n133 dd_02.n118 26.6872
R1109 dd_02.n93 dd_02.n33 26.345
R1110 dd_02.n178 dd_02.n156 18.0711
R1111 dd_02.n35 dd_02.n34 9.3005
R1112 dd_02.n34 dd_02.n33 9.3005
R1113 dd_02.n148 dd_02.n147 9.3005
R1114 dd_02.n147 dd_02.n146 9.3005
R1115 dd_02.n112 dd_02.n110 9.3005
R1116 dd_02.n112 dd_02.n111 9.3005
R1117 dd_02.n116 dd_02.n115 9.3005
R1118 dd_02.n117 dd_02.n116 9.3005
R1119 dd_02.n98 ring_100mV_0.mdls_inv_8.DD 7.37677
R1120 ring_100mV_0.mdls_inv_6.DD dd_02.n59 7.37677
R1121 ring_100mV_0.mdls_inv_4.DD dd_02.n46 7.37677
R1122 dd_02.n136 ring_100mV_0.mdls_inv_1.DD 7.37677
R1123 dd_02.n118 dd_02.n117 5.93087
R1124 dd_02.n46 ring_100mV_0.mdls_inv_5.DD 3.25474
R1125 dd_02.n59 ring_100mV_0.mdls_inv_7.DD 3.25474
R1126 ring_100mV_0.mdls_inv_9.DD dd_02.n98 3.25474
R1127 dd_02.n136 dd_02 3.25474
R1128 ring_100mV_0.DD dd_02 2.03619
R1129 dd_02.n166 dd_02.n156 1.95834
R1130 dd_02.n150 dd_02.n148 1.58284
R1131 dd_02.t2 dd_02.n89 1.255
R1132 dd_02.n115 dd_02.n113 1.10249
R1133 dd_02.t5 dd_02.n23 0.912865
R1134 ring_100mV_0.mdls_inv_3.DD dd_02.n35 0.848182
R1135 dd_02.n148 dd_02.n2 0.838796
R1136 dd_02.n114 dd_02.n1 0.765989
R1137 dd_02.n115 dd_02.n114 0.765989
R1138 dd_02.n173 dd_02.n166 0.753441
R1139 dd_02.n35 dd_02.n2 0.588624
R1140 dd_02.n180 dd_02.n151 0.518365
R1141 dd_02.n153 dd_02.n152 0.488
R1142 dd_02.n113 ring_100mV_0.mdls_inv_2.DD 0.226549
R1143 dd_02.n180 ring_100mV_0.ring_100mV_buffer_0.DD 0.204657
R1144 dd_02.n160 dd_02.n155 0.178278
R1145 ring_100mV_0.mdls_inv_2.DD dd_02.n112 0.14178
R1146 ring_100mV_0.DD dd_02.n180 0.130247
R1147 dd_02.n133 dd_02.t5 0.114546
R1148 dd_02.n93 dd_02.t2 0.114546
R1149 dd_02.n39 dd_02.n38 0.086406
R1150 dd_02.n129 dd_02.n128 0.086406
R1151 dd_02.n126 dd_02.n125 0.086406
R1152 dd_02.n123 dd_02.n122 0.086406
R1153 dd_02.n120 dd_02.n119 0.086406
R1154 dd_02.n68 dd_02.n67 0.086406
R1155 dd_02.n65 dd_02.n64 0.086406
R1156 dd_02.n52 dd_02.n51 0.086406
R1157 dd_02.n91 dd_02.n90 0.086406
R1158 dd_02.n25 dd_02.n24 0.086406
R1159 dd_02.n150 dd_02.n1 0.0570121
R1160 ring_100mV_0.ring_100mV_buffer_0.DD dd_02.n179 0.0290598
R1161 dd_02.n88 dd_02.n87 0.0204849
R1162 dd_02.n89 dd_02.n88 0.0204849
R1163 dd_02.n22 dd_02.n21 0.0202544
R1164 dd_02.n23 dd_02.n22 0.0202544
R1165 dd_02.n37 dd_02.n36 0.0194239
R1166 dd_02.n93 dd_02.n37 0.0194239
R1167 dd_02.n132 dd_02.n131 0.0194239
R1168 dd_02.n133 dd_02.n132 0.0194239
R1169 dd_02.n110 dd_02.n109 0.0183571
R1170 dd_02.n109 dd_02.n108 0.0165714
R1171 dd_02.n50 dd_02.n49 0.00996195
R1172 dd_02.n93 dd_02.n50 0.00996195
R1173 dd_02.n63 dd_02.n62 0.00996195
R1174 dd_02.n93 dd_02.n63 0.00996195
R1175 dd_02.n95 dd_02.n94 0.00996195
R1176 dd_02.n94 dd_02.n93 0.00996195
R1177 dd_02.n121 dd_02.n120 0.00996195
R1178 dd_02.n133 dd_02.n121 0.00996195
R1179 dd_02.n135 dd_02.n134 0.00996195
R1180 dd_02.n134 dd_02.n133 0.00996195
R1181 dd_02.n69 dd_02.n68 0.00996195
R1182 dd_02.n93 dd_02.n69 0.00996195
R1183 dd_02.n124 dd_02.n123 0.00996195
R1184 dd_02.n133 dd_02.n124 0.00996195
R1185 dd_02.n100 dd_02.n99 0.00996195
R1186 dd_02.n133 dd_02.n100 0.00996195
R1187 dd_02.n66 dd_02.n65 0.00996195
R1188 dd_02.n93 dd_02.n66 0.00996195
R1189 dd_02.n127 dd_02.n126 0.00996195
R1190 dd_02.n133 dd_02.n127 0.00996195
R1191 dd_02.n56 dd_02.n28 0.00996195
R1192 dd_02.n133 dd_02.n28 0.00996195
R1193 dd_02.n53 dd_02.n52 0.00996195
R1194 dd_02.n93 dd_02.n53 0.00996195
R1195 dd_02.n130 dd_02.n129 0.00996195
R1196 dd_02.n133 dd_02.n130 0.00996195
R1197 dd_02.n43 dd_02.n27 0.00996195
R1198 dd_02.n133 dd_02.n27 0.00996195
R1199 dd_02.n40 dd_02.n39 0.00996195
R1200 dd_02.n93 dd_02.n40 0.00996195
R1201 dd_02.n92 dd_02.n91 0.00996195
R1202 dd_02.n93 dd_02.n92 0.00996195
R1203 dd_02.n93 dd_02.n73 0.00996195
R1204 dd_02.n73 dd_02.n72 0.00996195
R1205 dd_02.n26 dd_02.n25 0.00996195
R1206 dd_02.n133 dd_02.n26 0.00996195
R1207 dd_02.n107 dd_02.n106 0.00705675
R1208 dd_02.n145 dd_02.n144 0.00705675
R1209 dd_02.n171 dd_02.n170 0.00696085
R1210 dd_02.n174 dd_02.n173 0.00696085
R1211 dd_02.n175 dd_02.n174 0.00696085
R1212 dd_02.n107 dd_02.n105 0.00693909
R1213 dd_02.n145 dd_02.n141 0.00693909
R1214 dd_02.n144 dd_02.n143 0.00655822
R1215 dd_02.n141 dd_02.n140 0.00644053
R1216 dd_02.n178 dd_02.n177 0.0063511
R1217 dd_02.n177 dd_02.n176 0.0063511
R1218 dd_02.n162 dd_02.n161 0.0063511
R1219 dd_02.n172 dd_02.n165 0.0046933
R1220 dd_02.n169 dd_02.n165 0.0046933
R1221 dd_02.n169 dd_02.n164 0.0046933
R1222 dd_02.n168 dd_02.n164 0.0046933
R1223 dd_02.n151 dd_02.n0 0.00407143
R1224 dd_02.n9 dd_02.n8 0.00347027
R1225 dd_02.n18 dd_02.n9 0.00347027
R1226 dd_02.n77 dd_02.n76 0.00347027
R1227 dd_02.n84 dd_02.n77 0.00347027
R1228 dd_02.n11 dd_02.n10 0.00347027
R1229 dd_02.n18 dd_02.n11 0.00347027
R1230 dd_02.n79 dd_02.n78 0.00347027
R1231 dd_02.n84 dd_02.n79 0.00347027
R1232 dd_02.n13 dd_02.n12 0.00347027
R1233 dd_02.n18 dd_02.n13 0.00347027
R1234 dd_02.n81 dd_02.n80 0.00347027
R1235 dd_02.n84 dd_02.n81 0.00347027
R1236 dd_02.n15 dd_02.n14 0.00347027
R1237 dd_02.n18 dd_02.n15 0.00347027
R1238 dd_02.n83 dd_02.n82 0.00347027
R1239 dd_02.n84 dd_02.n83 0.00347027
R1240 dd_02.n75 dd_02.n74 0.00347027
R1241 dd_02.n84 dd_02.n75 0.00347027
R1242 dd_02.n139 dd_02.n138 0.00347027
R1243 dd_02.n146 dd_02.n139 0.00347027
R1244 dd_02.n117 dd_02.n104 0.00347027
R1245 dd_02.n97 dd_02.n5 0.00347027
R1246 dd_02.n146 dd_02.n5 0.00347027
R1247 dd_02.n117 dd_02.n103 0.00347027
R1248 dd_02.n58 dd_02.n4 0.00347027
R1249 dd_02.n146 dd_02.n4 0.00347027
R1250 dd_02.n117 dd_02.n102 0.00347027
R1251 dd_02.n45 dd_02.n3 0.00347027
R1252 dd_02.n146 dd_02.n3 0.00347027
R1253 dd_02.n117 dd_02.n101 0.00347027
R1254 dd_02.n17 dd_02.n16 0.00347027
R1255 dd_02.n18 dd_02.n17 0.00347027
R1256 dd_02.n110 dd_02.n1 0.00335189
R1257 dd_02.n154 dd_02.n153 0.00314085
R1258 dd_02.n159 dd_02.n157 0.00294547
R1259 dd_02.n163 dd_02.n157 0.00294547
R1260 dd_02.n160 dd_02.n158 0.00294547
R1261 dd_02.n163 dd_02.n158 0.00294547
R1262 dd_02.n146 dd_02.n145 0.00100073
R1263 dd_02.n117 dd_02.n107 0.00100073
R1264 dd_02.n155 dd_02.n154 0.000500742
R1265 dd_02.n151 dd_02.n150 0.000500464
R1266 dd_02.n150 dd_02.n149 0.000500345
R1267 a_9754_13622.n4 a_9754_13622.t2 260.2
R1268 a_9754_13622.n2 a_9754_13622.t6 252.136
R1269 a_9754_13622.n0 a_9754_13622.t3 251.333
R1270 a_9754_13622.n3 a_9754_13622.n2 164.748
R1271 a_9754_13622.n0 a_9754_13622.t1 157.893
R1272 a_9754_13622.n1 a_9754_13622.t4 155.667
R1273 a_9754_13622.t5 a_9754_13622.n4 149.827
R1274 a_9754_13622.n3 a_9754_13622.n1 72.9605
R1275 a_9754_13622.n4 a_9754_13622.n3 9.14336
R1276 a_9754_13622.n1 a_9754_13622.n0 8.74717
R1277 a_9754_13622.n2 a_9754_13622.t0 3.16453
R1278 ldo_iref.n8 ldo_iref.t7 206.963
R1279 ldo_iref.n4 ldo_iref.t5 206.963
R1280 ldo_iref.n4 ldo_iref.t8 206.321
R1281 ldo_iref.n5 ldo_iref.t9 206.321
R1282 ldo_iref.n6 ldo_iref.t0 206.321
R1283 ldo_iref.n8 ldo_iref.t6 206.321
R1284 ldo_iref.n10 ldo_iref.t4 206.321
R1285 ldo_iref.n12 ldo_iref.t2 206.321
R1286 ldo_iref.t8 ldo_iref.n3 206.317
R1287 ldo_iref.t9 ldo_iref.n2 206.317
R1288 ldo_iref.t0 ldo_iref.n1 206.317
R1289 ldo_iref.t6 ldo_iref.n7 206.317
R1290 ldo_iref.t4 ldo_iref.n9 206.317
R1291 ldo_iref.t2 ldo_iref.n11 206.317
R1292 ldo_iref.n0 ldo_iref.t1 3.41293
R1293 ldo_iref.n0 ldo_iref.t3 3.41293
R1294 ldo_iref.n13 ldo_iref 1.7772
R1295 ldo_iref.n12 ldo_iref.n10 0.642396
R1296 ldo_iref.n10 ldo_iref.n8 0.642396
R1297 ldo_iref.n5 ldo_iref.n4 0.642396
R1298 ldo_iref.n6 ldo_iref.n5 0.642396
R1299 ldo_iref ldo_iref.n13 0.235123
R1300 ldo_iref.n13 ldo_iref.n6 0.192876
R1301 ldo_iref ldo_iref.n0 0.184094
R1302 ldo_iref.n13 ldo_iref.n12 0.183948
R1303 ring_100mV_0.mdls_inv_6.IN.n17 ring_100mV_0.mdls_inv_6.IN.t3 265.382
R1304 ring_100mV_0.mdls_inv_6.IN.n19 ring_100mV_0.mdls_inv_6.IN.n18 262.217
R1305 ring_100mV_0.mdls_inv_6.IN.n7 ring_100mV_0.mdls_inv_6.IN.t10 183.099
R1306 ring_100mV_0.mdls_inv_6.IN.n6 ring_100mV_0.mdls_inv_6.IN.t6 183.099
R1307 ring_100mV_0.mdls_inv_6.IN.t6 ring_100mV_0.mdls_inv_6.IN.n5 183.099
R1308 ring_100mV_0.mdls_inv_6.IN.n2 ring_100mV_0.mdls_inv_6.IN.t11 182.653
R1309 ring_100mV_0.mdls_inv_6.IN.t10 ring_100mV_0.mdls_inv_6.IN.n0 182.297
R1310 ring_100mV_0.mdls_inv_6.IN.n2 ring_100mV_0.mdls_inv_6.IN.t7 182.288
R1311 ring_100mV_0.mdls_inv_6.IN.n1 ring_100mV_0.mdls_inv_6.IN.t14 182.285
R1312 ring_100mV_0.mdls_inv_6.IN.n6 ring_100mV_0.mdls_inv_6.IN.t12 182.263
R1313 ring_100mV_0.mdls_inv_6.IN.t14 ring_100mV_0.mdls_inv_6.IN.n7 182.263
R1314 ring_100mV_0.mdls_inv_6.IN.t12 ring_100mV_0.mdls_inv_6.IN.n5 182.263
R1315 ring_100mV_0.mdls_inv_6.IN.n18 ring_100mV_0.mdls_inv_6.IN.t2 155.667
R1316 ring_100mV_0.mdls_inv_6.IN.n17 ring_100mV_0.mdls_inv_6.IN.t1 155.667
R1317 ring_100mV_0.mdls_inv_6.IN.t13 ring_100mV_0.mdls_inv_6.IN.n4 146.282
R1318 ring_100mV_0.mdls_inv_6.IN ring_100mV_0.mdls_inv_6.IN.t9 145.889
R1319 ring_100mV_0.mdls_inv_6.IN.t9 ring_100mV_0.mdls_inv_6.IN.n10 145.857
R1320 ring_100mV_0.mdls_inv_6.IN.n8 ring_100mV_0.mdls_inv_6.IN.t13 145.851
R1321 ring_100mV_0.mdls_inv_6.IN.n12 ring_100mV_0.mdls_inv_6.IN.t5 135.911
R1322 ring_100mV_0.mdls_inv_6.IN.n15 ring_100mV_0.mdls_inv_6.IN.n14 122.928
R1323 ring_100mV_0.mdls_inv_6.IN.n18 ring_100mV_0.mdls_inv_6.IN.n17 109.715
R1324 ring_100mV_0.mdls_inv_6.IN.t15 ring_100mV_0.mdls_inv_6.IN.n13 98.2234
R1325 ring_100mV_0.mdls_inv_6.IN.n15 ring_100mV_0.mdls_inv_6.IN.t15 49.4098
R1326 ring_100mV_0.mdls_inv_6.IN.n3 ring_100mV_0.mdls_inv_6.IN.t8 45.8204
R1327 ring_100mV_0.mdls_inv_6.IN.n12 ring_100mV_0.mdls_inv_6.IN.n3 28.5785
R1328 ring_100mV_0.mdls_inv_6.IN.n14 ring_100mV_0.mdls_inv_6.IN.t0 28.5685
R1329 ring_100mV_0.mdls_inv_6.IN.t5 ring_100mV_0.mdls_inv_6.IN.n11 19.7637
R1330 ring_100mV_0.mdls_inv_6.IN.n16 ring_100mV_0.mdls_inv_6.IN.n15 5.00095
R1331 ring_100mV_0.mdls_inv_6.IN.n9 ring_100mV_0.mdls_inv_6.IN.n4 4.13208
R1332 ring_100mV_0.mdls_inv_6.IN.n19 ring_100mV_0.mdls_inv_6.IN.t4 3.16453
R1333 ring_100mV_0.mdls_inv_6.IN.n16 ring_100mV_0.mdls_inv_6.IN.n2 1.3453
R1334 ring_100mV_0.mdls_inv_8.OUT ring_100mV_0.mdls_inv_6.IN.n19 1.29092
R1335 ring_100mV_0.mdls_inv_6.IN.n13 ring_100mV_0.mdls_inv_6.IN.n12 1.06388
R1336 ring_100mV_0.mdls_inv_6.IN.n7 ring_100mV_0.mdls_inv_6.IN.n6 0.835457
R1337 ring_100mV_0.mdls_inv_6.IN.n1 ring_100mV_0.mdls_inv_6.IN.n5 0.813812
R1338 ring_100mV_0.mdls_inv_6.IN.n1 ring_100mV_0.mdls_inv_6.IN.n0 0.810242
R1339 ring_100mV_0.mdls_inv_6.IN.n10 ring_100mV_0.mdls_inv_6.IN.n9 0.607643
R1340 ring_100mV_0.mdls_inv_6.IN ring_100mV_0.mdls_inv_6.IN.n4 0.454134
R1341 ring_100mV_0.mdls_inv_6.IN.n9 ring_100mV_0.mdls_inv_6.IN.n8 0.43198
R1342 ring_100mV_0.mdls_inv_6.IN.n11 ring_100mV_0.mdls_inv_6.IN 0.339159
R1343 ring_100mV_0.mdls_inv_6.IN.n8 ring_100mV_0.mdls_inv_6.IN.n1 0.320167
R1344 ring_100mV_0.mdls_inv_6.IN.n10 ring_100mV_0.mdls_inv_6.IN.n0 0.21421
R1345 ring_100mV_0.mdls_inv_8.OUT ring_100mV_0.mdls_inv_6.IN.n16 0.184521
R1346 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n0 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t4 21.4396
R1347 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n0 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t6 18.8004
R1348 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n1 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t5 18.8004
R1349 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n2 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t3 18.8004
R1350 iref_2nA_0.iref_2nA_mirrors_0.Ip1 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t2 11.5886
R1351 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n3 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t0 11.5885
R1352 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n4 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t1 8.4133
R1353 iref_2nA_0.iref_2nA_mirrors_0.Ip1 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n2 7.65117
R1354 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n3 iref_2nA_0.iref_2nA_mirrors_0.Ip1 3.82182
R1355 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n1 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n0 2.63976
R1356 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n2 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n1 2.63976
R1357 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n4 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n3 1.93205
R1358 iref_2nA_0.iref_2nA_igenerator_0.Ip1 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n4 0.573
R1359 ring_100mV_0.mdls_inv_3.OUT.n17 ring_100mV_0.mdls_inv_3.OUT.n9 368.413
R1360 ring_100mV_0.mdls_inv_3.OUT.n22 ring_100mV_0.mdls_inv_3.OUT.t0 265.382
R1361 ring_100mV_0.mdls_inv_3.OUT.n24 ring_100mV_0.mdls_inv_3.OUT.n23 262.217
R1362 ring_100mV_0.mdls_inv_3.OUT.n10 ring_100mV_0.mdls_inv_3.OUT.t14 251.451
R1363 ring_100mV_0.mdls_inv_3.OUT.n1 ring_100mV_0.mdls_inv_3.OUT.t5 182.653
R1364 ring_100mV_0.mdls_inv_3.OUT.n1 ring_100mV_0.mdls_inv_3.OUT.t10 182.288
R1365 ring_100mV_0.mdls_inv_3.OUT.n10 ring_100mV_0.mdls_inv_3.OUT.t9 182.262
R1366 ring_100mV_0.mdls_inv_3.OUT.n11 ring_100mV_0.mdls_inv_3.OUT.t16 182.262
R1367 ring_100mV_0.mdls_inv_3.OUT.n12 ring_100mV_0.mdls_inv_3.OUT.t12 182.262
R1368 ring_100mV_0.mdls_inv_3.OUT.n13 ring_100mV_0.mdls_inv_3.OUT.t17 182.262
R1369 ring_100mV_0.mdls_inv_3.OUT.n14 ring_100mV_0.mdls_inv_3.OUT.t13 182.262
R1370 ring_100mV_0.mdls_inv_3.OUT.n15 ring_100mV_0.mdls_inv_3.OUT.t8 182.262
R1371 ring_100mV_0.mdls_inv_3.OUT.n16 ring_100mV_0.mdls_inv_3.OUT.t15 182.262
R1372 ring_100mV_0.mdls_inv_3.OUT.n23 ring_100mV_0.mdls_inv_3.OUT.t2 155.667
R1373 ring_100mV_0.mdls_inv_3.OUT.n22 ring_100mV_0.mdls_inv_3.OUT.t4 155.667
R1374 ring_100mV_0.mdls_inv_3.OUT.n20 ring_100mV_0.mdls_inv_3.OUT.n19 122.928
R1375 ring_100mV_0.mdls_inv_3.OUT.n23 ring_100mV_0.mdls_inv_3.OUT.n22 109.715
R1376 ring_100mV_0.mdls_inv_3.OUT.t7 ring_100mV_0.mdls_inv_3.OUT.n18 98.2234
R1377 ring_100mV_0.mdls_inv_3.OUT.n9 ring_100mV_0.mdls_inv_3.OUT.n8 72.1132
R1378 ring_100mV_0.mdls_inv_3.OUT.n8 ring_100mV_0.mdls_inv_3.OUT.n7 72.1132
R1379 ring_100mV_0.mdls_inv_3.OUT.n7 ring_100mV_0.mdls_inv_3.OUT.n6 72.1132
R1380 ring_100mV_0.mdls_inv_3.OUT.n6 ring_100mV_0.mdls_inv_3.OUT.n5 72.1132
R1381 ring_100mV_0.mdls_inv_3.OUT.n5 ring_100mV_0.mdls_inv_3.OUT.n4 72.1132
R1382 ring_100mV_0.mdls_inv_3.OUT.n4 ring_100mV_0.mdls_inv_3.OUT.n3 72.1132
R1383 ring_100mV_0.mdls_inv_3.OUT.n16 ring_100mV_0.mdls_inv_3.OUT.n15 69.1897
R1384 ring_100mV_0.mdls_inv_3.OUT.n15 ring_100mV_0.mdls_inv_3.OUT.n14 69.1897
R1385 ring_100mV_0.mdls_inv_3.OUT.n14 ring_100mV_0.mdls_inv_3.OUT.n13 69.1897
R1386 ring_100mV_0.mdls_inv_3.OUT.n13 ring_100mV_0.mdls_inv_3.OUT.n12 69.1897
R1387 ring_100mV_0.mdls_inv_3.OUT.n12 ring_100mV_0.mdls_inv_3.OUT.n11 69.1897
R1388 ring_100mV_0.mdls_inv_3.OUT.n11 ring_100mV_0.mdls_inv_3.OUT.n10 69.1897
R1389 ring_100mV_0.mdls_inv_3.OUT.n17 ring_100mV_0.mdls_inv_3.OUT.n16 62.0129
R1390 ring_100mV_0.mdls_inv_3.OUT.n20 ring_100mV_0.mdls_inv_3.OUT.t7 49.4098
R1391 ring_100mV_0.mdls_inv_3.OUT.n2 ring_100mV_0.mdls_inv_3.OUT.t6 36.7438
R1392 ring_100mV_0.mdls_inv_3.OUT.n2 ring_100mV_0.mdls_inv_3.OUT.t11 32.5647
R1393 ring_100mV_0.mdls_inv_3.OUT.n19 ring_100mV_0.mdls_inv_3.OUT.t3 28.5685
R1394 ring_100mV_0.mdls_inv_3.OUT.n0 ring_100mV_0.mdls_inv_3.OUT.n17 27.9962
R1395 ring_100mV_0.mdls_inv_3.OUT.n0 ring_100mV_0.mdls_inv_3.OUT.n2 6.45024
R1396 ring_100mV_0.mdls_inv_3.OUT.n21 ring_100mV_0.mdls_inv_3.OUT.n20 5.00095
R1397 ring_100mV_0.mdls_inv_3.OUT.n24 ring_100mV_0.mdls_inv_3.OUT.t1 3.16453
R1398 ring_100mV_0.mdls_inv_3.OUT.n18 ring_100mV_0.mdls_inv_3.OUT.n0 2.08823
R1399 ring_100mV_0.mdls_inv_3.OUT.n21 ring_100mV_0.mdls_inv_3.OUT.n1 1.3453
R1400 ring_100mV_0.mdls_inv_3.OUT ring_100mV_0.mdls_inv_3.OUT.n24 1.29092
R1401 ring_100mV_0.mdls_inv_3.OUT ring_100mV_0.mdls_inv_3.OUT.n21 0.184521
R1402 ring_100mV_0.mdls_inv_3.OUT.n0 ring_100mV_0.ring_100mV_buffer_0.IN 0.156641
R1403 a_16150_16902.n7 a_16150_16902.t4 177.476
R1404 a_16150_16902.n6 a_16150_16902.t2 177.371
R1405 a_16150_16902.n5 a_16150_16902.t6 31.4497
R1406 a_16150_16902.n0 a_16150_16902.t0 17.6491
R1407 a_16150_16902.n3 a_16150_16902.t1 10.2714
R1408 a_16150_16902.t5 a_16150_16902.n7 4.93845
R1409 a_16150_16902.n0 a_16150_16902.t3 2.90106
R1410 a_16150_16902.n5 a_16150_16902.n0 0.941548
R1411 a_16150_16902.n3 a_16150_16902.n2 0.923627
R1412 a_16150_16902.n0 a_16150_16902.n4 0.836115
R1413 a_16150_16902.n4 a_16150_16902.n1 0.773938
R1414 a_16150_16902.n6 a_16150_16902.n5 0.288679
R1415 a_16150_16902.n4 a_16150_16902.n3 0.224162
R1416 a_16150_16902.n7 a_16150_16902.n6 0.0975343
R1417 vref.n0 vref.t0 636.341
R1418 vref.n3 vref.n0 365.553
R1419 vref.n2 vref.n1 365.553
R1420 vref.n3 vref.n2 365.553
R1421 vref.n4 vref.t3 21.3068
R1422 vref.n6 vref.n5 11.9344
R1423 vref.n4 vref.t4 10.1983
R1424 vref.n3 vref.t1 3.32227
R1425 vref.n1 vref.t2 3.32227
R1426 vref.n6 vref.n3 2.59757
R1427 vref.n5 vref.n4 1.60834
R1428 vref.n5 vref 0.829256
R1429 vref vref.n6 0.0165714
R1430 a_14834_9380.n0 a_14834_9380.t2 7.40825
R1431 a_14834_9380.n0 a_14834_9380.t3 4.70699
R1432 a_14834_9380.t6 a_14834_9380.n5 4.53569
R1433 a_14834_9380.n2 a_14834_9380.t5 4.53369
R1434 a_14834_9380.n3 a_14834_9380.t4 4.38957
R1435 a_14834_9380.n4 a_14834_9380.t7 4.3873
R1436 a_14834_9380.n1 a_14834_9380.t1 4.26166
R1437 a_14834_9380.n1 a_14834_9380.t0 4.06962
R1438 a_14834_9380.n4 a_14834_9380.n3 2.26478
R1439 a_14834_9380.n2 a_14834_9380.n1 2.0915
R1440 a_14834_9380.n5 a_14834_9380.n0 0.66715
R1441 a_14834_9380.n3 a_14834_9380.n2 0.1505
R1442 a_14834_9380.n5 a_14834_9380.n4 0.144506
R1443 a_9754_8624.n2 a_9754_8624.t6 260.2
R1444 a_9754_8624.n4 a_9754_8624.t0 252.136
R1445 a_9754_8624.n0 a_9754_8624.t2 251.333
R1446 a_9754_8624.n4 a_9754_8624.n3 164.748
R1447 a_9754_8624.n0 a_9754_8624.t3 157.893
R1448 a_9754_8624.n1 a_9754_8624.t1 155.667
R1449 a_9754_8624.n2 a_9754_8624.t5 149.827
R1450 a_9754_8624.n3 a_9754_8624.n1 72.9605
R1451 a_9754_8624.n3 a_9754_8624.n2 9.14336
R1452 a_9754_8624.n1 a_9754_8624.n0 8.74717
R1453 a_9754_8624.t4 a_9754_8624.n4 3.16453
R1454 ring_100mV_0.mdls_inv_0.OUT.n0 ring_100mV_0.mdls_inv_0.OUT.t2 265.382
R1455 ring_100mV_0.mdls_inv_0.OUT.n2 ring_100mV_0.mdls_inv_0.OUT.n1 262.217
R1456 ring_100mV_0.mdls_inv_0.OUT.n9 ring_100mV_0.mdls_inv_0.OUT.t7 183.099
R1457 ring_100mV_0.mdls_inv_0.OUT.n8 ring_100mV_0.mdls_inv_0.OUT.t12 183.099
R1458 ring_100mV_0.mdls_inv_0.OUT.t12 ring_100mV_0.mdls_inv_0.OUT.n7 183.099
R1459 ring_100mV_0.mdls_inv_0.OUT.n3 ring_100mV_0.mdls_inv_0.OUT.t15 182.653
R1460 ring_100mV_0.mdls_inv_0.OUT.t7 ring_100mV_0.mdls_inv_0.OUT.n6 182.297
R1461 ring_100mV_0.mdls_inv_0.OUT.n3 ring_100mV_0.mdls_inv_0.OUT.t9 182.288
R1462 ring_100mV_0.mdls_inv_0.OUT.n10 ring_100mV_0.mdls_inv_0.OUT.t6 182.285
R1463 ring_100mV_0.mdls_inv_0.OUT.n8 ring_100mV_0.mdls_inv_0.OUT.t13 182.263
R1464 ring_100mV_0.mdls_inv_0.OUT.t6 ring_100mV_0.mdls_inv_0.OUT.n9 182.263
R1465 ring_100mV_0.mdls_inv_0.OUT.t13 ring_100mV_0.mdls_inv_0.OUT.n7 182.263
R1466 ring_100mV_0.mdls_inv_0.OUT.n1 ring_100mV_0.mdls_inv_0.OUT.t0 155.667
R1467 ring_100mV_0.mdls_inv_0.OUT.n0 ring_100mV_0.mdls_inv_0.OUT.t3 155.667
R1468 ring_100mV_0.mdls_inv_0.OUT.t8 ring_100mV_0.mdls_inv_0.OUT.n5 146.282
R1469 ring_100mV_0.mdls_inv_0.OUT.n15 ring_100mV_0.mdls_inv_0.OUT.t14 145.889
R1470 ring_100mV_0.mdls_inv_0.OUT.t14 ring_100mV_0.mdls_inv_0.OUT.n14 145.857
R1471 ring_100mV_0.mdls_inv_0.OUT.n12 ring_100mV_0.mdls_inv_0.OUT.t8 145.851
R1472 ring_100mV_0.mdls_inv_0.OUT.n17 ring_100mV_0.mdls_inv_0.OUT.t11 135.911
R1473 ring_100mV_0.mdls_inv_0.OUT.n20 ring_100mV_0.mdls_inv_0.OUT.n19 122.928
R1474 ring_100mV_0.mdls_inv_0.OUT.n1 ring_100mV_0.mdls_inv_0.OUT.n0 109.715
R1475 ring_100mV_0.mdls_inv_0.OUT.t10 ring_100mV_0.mdls_inv_0.OUT.n18 98.2234
R1476 ring_100mV_0.mdls_inv_0.OUT.n20 ring_100mV_0.mdls_inv_0.OUT.t10 49.4098
R1477 ring_100mV_0.mdls_inv_0.OUT.n4 ring_100mV_0.mdls_inv_0.OUT.t5 45.8204
R1478 ring_100mV_0.mdls_inv_0.OUT.n17 ring_100mV_0.mdls_inv_0.OUT.n4 28.5785
R1479 ring_100mV_0.mdls_inv_0.OUT.n19 ring_100mV_0.mdls_inv_0.OUT.t4 28.5685
R1480 ring_100mV_0.mdls_inv_0.OUT.t11 ring_100mV_0.mdls_inv_0.OUT.n16 19.7637
R1481 ring_100mV_0.mdls_inv_0.OUT.n18 ring_100mV_0.mdls_inv_0.OUT.n17 5.198
R1482 ring_100mV_0.mdls_inv_0.OUT.n21 ring_100mV_0.mdls_inv_0.OUT.n20 5.00095
R1483 ring_100mV_0.mdls_inv_0.OUT.n13 ring_100mV_0.mdls_inv_0.OUT.n5 4.13208
R1484 ring_100mV_0.mdls_inv_0.OUT.n2 ring_100mV_0.mdls_inv_0.OUT.t1 3.16453
R1485 ring_100mV_0.mdls_inv_0.OUT ring_100mV_0.mdls_inv_0.OUT.n2 1.36143
R1486 ring_100mV_0.mdls_inv_0.OUT.n21 ring_100mV_0.mdls_inv_0.OUT.n3 1.34518
R1487 ring_100mV_0.mdls_inv_0.OUT.n9 ring_100mV_0.mdls_inv_0.OUT.n8 0.835457
R1488 ring_100mV_0.mdls_inv_0.OUT.n11 ring_100mV_0.mdls_inv_0.OUT.n7 0.813812
R1489 ring_100mV_0.mdls_inv_0.OUT.n10 ring_100mV_0.mdls_inv_0.OUT.n6 0.810242
R1490 ring_100mV_0.mdls_inv_0.OUT.n14 ring_100mV_0.mdls_inv_0.OUT.n13 0.607643
R1491 ring_100mV_0.mdls_inv_0.OUT.n13 ring_100mV_0.mdls_inv_0.OUT.n12 0.43198
R1492 ring_100mV_0.mdls_inv_0.OUT.n16 ring_100mV_0.mdls_inv_1.IN 0.339159
R1493 ring_100mV_0.mdls_inv_0.OUT.n15 ring_100mV_0.mdls_inv_0.OUT.n5 0.333833
R1494 ring_100mV_0.mdls_inv_0.OUT.n12 ring_100mV_0.mdls_inv_0.OUT.n11 0.21421
R1495 ring_100mV_0.mdls_inv_0.OUT.n14 ring_100mV_0.mdls_inv_0.OUT.n6 0.21421
R1496 ring_100mV_0.mdls_inv_1.IN ring_100mV_0.mdls_inv_0.OUT.n15 0.120801
R1497 ring_100mV_0.mdls_inv_0.OUT ring_100mV_0.mdls_inv_0.OUT.n21 0.114008
R1498 ring_100mV_0.mdls_inv_0.OUT.n11 ring_100mV_0.mdls_inv_0.OUT.n10 0.106457
R1499 ring_100mV_0.mdls_inv_1.OUT.n17 ring_100mV_0.mdls_inv_1.OUT.t3 265.382
R1500 ring_100mV_0.mdls_inv_1.OUT.n19 ring_100mV_0.mdls_inv_1.OUT.n18 262.217
R1501 ring_100mV_0.mdls_inv_1.OUT.n7 ring_100mV_0.mdls_inv_1.OUT.t5 183.099
R1502 ring_100mV_0.mdls_inv_1.OUT.n6 ring_100mV_0.mdls_inv_1.OUT.t11 183.099
R1503 ring_100mV_0.mdls_inv_1.OUT.t11 ring_100mV_0.mdls_inv_1.OUT.n5 183.099
R1504 ring_100mV_0.mdls_inv_1.OUT.n2 ring_100mV_0.mdls_inv_1.OUT.t9 182.653
R1505 ring_100mV_0.mdls_inv_1.OUT.t5 ring_100mV_0.mdls_inv_1.OUT.n0 182.297
R1506 ring_100mV_0.mdls_inv_1.OUT.n2 ring_100mV_0.mdls_inv_1.OUT.t15 182.288
R1507 ring_100mV_0.mdls_inv_1.OUT.n1 ring_100mV_0.mdls_inv_1.OUT.t7 182.285
R1508 ring_100mV_0.mdls_inv_1.OUT.n6 ring_100mV_0.mdls_inv_1.OUT.t8 182.263
R1509 ring_100mV_0.mdls_inv_1.OUT.t7 ring_100mV_0.mdls_inv_1.OUT.n7 182.263
R1510 ring_100mV_0.mdls_inv_1.OUT.t8 ring_100mV_0.mdls_inv_1.OUT.n5 182.263
R1511 ring_100mV_0.mdls_inv_1.OUT.n17 ring_100mV_0.mdls_inv_1.OUT.t4 155.667
R1512 ring_100mV_0.mdls_inv_1.OUT.n18 ring_100mV_0.mdls_inv_1.OUT.t0 155.667
R1513 ring_100mV_0.mdls_inv_1.OUT.t10 ring_100mV_0.mdls_inv_1.OUT.n4 146.282
R1514 ring_100mV_0.mdls_inv_8.IN ring_100mV_0.mdls_inv_1.OUT.t13 145.889
R1515 ring_100mV_0.mdls_inv_1.OUT.t13 ring_100mV_0.mdls_inv_1.OUT.n10 145.857
R1516 ring_100mV_0.mdls_inv_1.OUT.n8 ring_100mV_0.mdls_inv_1.OUT.t10 145.851
R1517 ring_100mV_0.mdls_inv_1.OUT.n12 ring_100mV_0.mdls_inv_1.OUT.t12 135.911
R1518 ring_100mV_0.mdls_inv_1.OUT.n15 ring_100mV_0.mdls_inv_1.OUT.n14 122.928
R1519 ring_100mV_0.mdls_inv_1.OUT.n18 ring_100mV_0.mdls_inv_1.OUT.n17 109.715
R1520 ring_100mV_0.mdls_inv_1.OUT.t14 ring_100mV_0.mdls_inv_1.OUT.n13 98.2234
R1521 ring_100mV_0.mdls_inv_1.OUT.n15 ring_100mV_0.mdls_inv_1.OUT.t14 49.4098
R1522 ring_100mV_0.mdls_inv_1.OUT.n3 ring_100mV_0.mdls_inv_1.OUT.t6 45.8204
R1523 ring_100mV_0.mdls_inv_1.OUT.n12 ring_100mV_0.mdls_inv_1.OUT.n3 28.5785
R1524 ring_100mV_0.mdls_inv_1.OUT.n14 ring_100mV_0.mdls_inv_1.OUT.t2 28.5685
R1525 ring_100mV_0.mdls_inv_1.OUT.t12 ring_100mV_0.mdls_inv_1.OUT.n11 19.7637
R1526 ring_100mV_0.mdls_inv_1.OUT.n16 ring_100mV_0.mdls_inv_1.OUT.n15 5.00095
R1527 ring_100mV_0.mdls_inv_1.OUT.n9 ring_100mV_0.mdls_inv_1.OUT.n4 4.13208
R1528 ring_100mV_0.mdls_inv_1.OUT.n19 ring_100mV_0.mdls_inv_1.OUT.t1 3.16453
R1529 ring_100mV_0.mdls_inv_1.OUT.n13 ring_100mV_0.mdls_inv_1.OUT.n12 2.84116
R1530 ring_100mV_0.mdls_inv_1.OUT.n16 ring_100mV_0.mdls_inv_1.OUT.n2 1.3453
R1531 ring_100mV_0.mdls_inv_1.OUT ring_100mV_0.mdls_inv_1.OUT.n19 1.29092
R1532 ring_100mV_0.mdls_inv_1.OUT.n7 ring_100mV_0.mdls_inv_1.OUT.n6 0.835457
R1533 ring_100mV_0.mdls_inv_1.OUT.n1 ring_100mV_0.mdls_inv_1.OUT.n5 0.813812
R1534 ring_100mV_0.mdls_inv_1.OUT.n1 ring_100mV_0.mdls_inv_1.OUT.n0 0.810242
R1535 ring_100mV_0.mdls_inv_1.OUT.n10 ring_100mV_0.mdls_inv_1.OUT.n9 0.607643
R1536 ring_100mV_0.mdls_inv_8.IN ring_100mV_0.mdls_inv_1.OUT.n4 0.454134
R1537 ring_100mV_0.mdls_inv_1.OUT.n9 ring_100mV_0.mdls_inv_1.OUT.n8 0.43198
R1538 ring_100mV_0.mdls_inv_1.OUT.n11 ring_100mV_0.mdls_inv_8.IN 0.339159
R1539 ring_100mV_0.mdls_inv_1.OUT.n8 ring_100mV_0.mdls_inv_1.OUT.n1 0.320167
R1540 ring_100mV_0.mdls_inv_1.OUT.n10 ring_100mV_0.mdls_inv_1.OUT.n0 0.21421
R1541 ring_100mV_0.mdls_inv_1.OUT ring_100mV_0.mdls_inv_1.OUT.n16 0.184521
R1542 a_15054_7578.n1 a_15054_7578.t3 32.4466
R1543 a_15054_7578.n0 a_15054_7578.t1 32.4466
R1544 a_15054_7578.t2 a_15054_7578.t7 19.1411
R1545 a_15054_7578.t0 a_15054_7578.t6 19.1411
R1546 a_15054_7578.n4 a_15054_7578.t4 10.1828
R1547 a_15054_7578.n3 a_15054_7578.t2 9.48031
R1548 a_15054_7578.n2 a_15054_7578.t0 9.48031
R1549 a_15054_7578.n4 a_15054_7578.n1 5.92365
R1550 a_15054_7578.t5 a_15054_7578.n4 5.36911
R1551 a_15054_7578.n0 a_15054_7578.n2 0.351043
R1552 a_15054_7578.n1 a_15054_7578.n3 0.351043
R1553 a_15054_7578.n1 a_15054_7578.n0 0.100294
R1554 a_14490_9380.n0 a_14490_9380.t4 191.636
R1555 a_14490_9380.n0 a_14490_9380.t0 34.661
R1556 a_14490_9380.n0 a_14490_9380.t1 33.291
R1557 a_14490_9380.t2 a_14490_9380.n1 4.51459
R1558 a_14490_9380.n1 a_14490_9380.t3 3.35375
R1559 a_14490_9380.t5 a_14490_9380.n0 2.51069
R1560 a_14490_9380.n1 a_14490_9380.t5 1.37236
R1561 a_5930_7513.n1 a_5930_7513.t1 260.2
R1562 a_5930_7513.n0 a_5930_7513.t6 252.136
R1563 a_5930_7513.n3 a_5930_7513.t2 251.333
R1564 a_5930_7513.n2 a_5930_7513.n0 164.748
R1565 a_5930_7513.n3 a_5930_7513.t4 157.893
R1566 a_5930_7513.t3 a_5930_7513.n4 155.667
R1567 a_5930_7513.n1 a_5930_7513.t0 149.827
R1568 a_5930_7513.n4 a_5930_7513.n2 72.9605
R1569 a_5930_7513.n2 a_5930_7513.n1 9.14336
R1570 a_5930_7513.n4 a_5930_7513.n3 8.74717
R1571 a_5930_7513.n0 a_5930_7513.t5 3.16453
R1572 a_9754_11956.n0 a_9754_11956.t1 260.2
R1573 a_9754_11956.n1 a_9754_11956.t0 252.136
R1574 a_9754_11956.t4 a_9754_11956.n4 251.333
R1575 a_9754_11956.n2 a_9754_11956.n1 164.748
R1576 a_9754_11956.n4 a_9754_11956.t5 157.893
R1577 a_9754_11956.n3 a_9754_11956.t2 155.667
R1578 a_9754_11956.n0 a_9754_11956.t3 149.827
R1579 a_9754_11956.n3 a_9754_11956.n2 72.9605
R1580 a_9754_11956.n2 a_9754_11956.n0 9.14336
R1581 a_9754_11956.n4 a_9754_11956.n3 8.74717
R1582 a_9754_11956.n1 a_9754_11956.t6 3.16453
R1583 a_955_10311.n0 a_955_10311.t1 57.4135
R1584 a_955_10311.n0 a_955_10311.t2 9.98238
R1585 a_955_10311.t0 a_955_10311.n0 9.18355
R1586 a_5712_16467.n26 a_5712_16467.t22 332.849
R1587 a_5712_16467.n6 a_5712_16467.n5 212.389
R1588 a_5712_16467.n6 a_5712_16467.t12 182.262
R1589 a_5712_16467.n7 a_5712_16467.t25 182.262
R1590 a_5712_16467.n8 a_5712_16467.t16 182.262
R1591 a_5712_16467.n9 a_5712_16467.t29 182.262
R1592 a_5712_16467.n10 a_5712_16467.t20 182.262
R1593 a_5712_16467.n17 a_5712_16467.t11 182.262
R1594 a_5712_16467.t11 a_5712_16467.n16 182.262
R1595 a_5712_16467.n18 a_5712_16467.t23 182.262
R1596 a_5712_16467.n21 a_5712_16467.t14 182.262
R1597 a_5712_16467.t14 a_5712_16467.n20 182.262
R1598 a_5712_16467.n22 a_5712_16467.t27 182.262
R1599 a_5712_16467.n25 a_5712_16467.t18 182.262
R1600 a_5712_16467.t18 a_5712_16467.n24 182.262
R1601 a_5712_16467.n33 a_5712_16467.t13 182.262
R1602 a_5712_16467.t13 a_5712_16467.n32 182.262
R1603 a_5712_16467.n28 a_5712_16467.t26 182.262
R1604 a_5712_16467.n27 a_5712_16467.t17 182.262
R1605 a_5712_16467.n26 a_5712_16467.t10 182.262
R1606 a_5712_16467.n30 a_5712_16467.n29 150.589
R1607 a_5712_16467.n31 a_5712_16467.n30 150.589
R1608 a_5712_16467.n32 a_5712_16467.n31 150.589
R1609 a_5712_16467.n24 a_5712_16467.n23 150.589
R1610 a_5712_16467.n20 a_5712_16467.n19 150.589
R1611 a_5712_16467.n16 a_5712_16467.n15 150.589
R1612 a_5712_16467.n15 a_5712_16467.n14 150.589
R1613 a_5712_16467.n14 a_5712_16467.n13 150.589
R1614 a_5712_16467.n13 a_5712_16467.n12 150.589
R1615 a_5712_16467.n12 a_5712_16467.n11 150.589
R1616 a_5712_16467.n25 a_5712_16467.n22 150.589
R1617 a_5712_16467.n22 a_5712_16467.n21 150.589
R1618 a_5712_16467.n21 a_5712_16467.n18 150.589
R1619 a_5712_16467.n18 a_5712_16467.n17 150.589
R1620 a_5712_16467.n17 a_5712_16467.n10 150.589
R1621 a_5712_16467.n10 a_5712_16467.n9 150.589
R1622 a_5712_16467.n9 a_5712_16467.n8 150.589
R1623 a_5712_16467.n8 a_5712_16467.n7 150.589
R1624 a_5712_16467.n7 a_5712_16467.n6 150.589
R1625 a_5712_16467.n27 a_5712_16467.n26 150.589
R1626 a_5712_16467.n28 a_5712_16467.n27 150.589
R1627 a_5712_16467.n33 a_5712_16467.n28 150.589
R1628 a_5712_16467.n37 a_5712_16467.n36 150.589
R1629 a_5712_16467.n39 a_5712_16467.n38 150.589
R1630 a_5712_16467.n36 a_5712_16467.n35 96.6009
R1631 a_5712_16467.n41 a_5712_16467.n40 87.4672
R1632 a_5712_16467.n41 a_5712_16467.n37 66.2593
R1633 a_5712_16467.n40 a_5712_16467.n39 66.2593
R1634 a_5712_16467.n42 a_5712_16467.n41 66.2593
R1635 a_5712_16467.n37 a_5712_16467.t15 49.4098
R1636 a_5712_16467.n36 a_5712_16467.t28 49.4098
R1637 a_5712_16467.n42 a_5712_16467.t24 49.4098
R1638 a_5712_16467.n34 a_5712_16467.n33 46.6829
R1639 a_5712_16467.n35 a_5712_16467.t19 42.6645
R1640 a_5712_16467.n5 a_5712_16467.t21 40.6427
R1641 a_5712_16467.n34 a_5712_16467.n25 38.777
R1642 a_5712_16467.n44 a_5712_16467.n34 32.5457
R1643 a_5712_16467.n44 a_5712_16467.t0 30.2238
R1644 a_5712_16467.n43 a_5712_16467.t1 28.5701
R1645 a_5712_16467.n0 a_5712_16467.t5 5.95384
R1646 a_5712_16467.n45 a_5712_16467.n44 4.84496
R1647 a_5712_16467.t9 a_5712_16467.n46 4.60076
R1648 a_5712_16467.n45 a_5712_16467.t4 4.60076
R1649 a_5712_16467.n0 a_5712_16467.t8 4.59778
R1650 a_5712_16467.n1 a_5712_16467.t3 4.59778
R1651 a_5712_16467.n2 a_5712_16467.t7 4.59778
R1652 a_5712_16467.n3 a_5712_16467.t2 4.59778
R1653 a_5712_16467.n4 a_5712_16467.t6 4.59778
R1654 a_5712_16467.n44 a_5712_16467.n43 2.10396
R1655 a_5712_16467.n43 a_5712_16467.n42 1.96379
R1656 a_5712_16467.n1 a_5712_16467.n0 1.35656
R1657 a_5712_16467.n2 a_5712_16467.n1 1.35656
R1658 a_5712_16467.n3 a_5712_16467.n2 1.35656
R1659 a_5712_16467.n4 a_5712_16467.n3 1.35656
R1660 a_5712_16467.n46 a_5712_16467.n4 1.33027
R1661 a_5712_16467.n46 a_5712_16467.n45 1.31668
R1662 ring_out.n0 ring_out.t1 30.4433
R1663 ring_out.n2 ring_out.t2 29.7591
R1664 ring_out.n0 ring_out.t3 29.2657
R1665 ring_out.n1 ring_out.t0 29.2657
R1666 ring_out.n3 ring_out.t10 5.86456
R1667 ring_out ring_out.t9 4.50884
R1668 ring_out.n3 ring_out.t17 4.5085
R1669 ring_out.n4 ring_out.t7 4.5085
R1670 ring_out.n5 ring_out.t14 4.5085
R1671 ring_out.n6 ring_out.t4 4.5085
R1672 ring_out.n7 ring_out.t11 4.5085
R1673 ring_out.n8 ring_out.t18 4.5085
R1674 ring_out.n9 ring_out.t8 4.5085
R1675 ring_out.n10 ring_out.t15 4.5085
R1676 ring_out.n11 ring_out.t5 4.5085
R1677 ring_out.n12 ring_out.t12 4.5085
R1678 ring_out.n13 ring_out.t16 4.5085
R1679 ring_out.n14 ring_out.t6 4.5085
R1680 ring_out.n16 ring_out.t19 4.4579
R1681 ring_out.n15 ring_out.t13 4.4579
R1682 ring_out.n1 ring_out.n0 2.18471
R1683 ring_out.n17 ring_out 2.0232
R1684 ring_out.n4 ring_out.n3 1.35656
R1685 ring_out.n5 ring_out.n4 1.35656
R1686 ring_out.n6 ring_out.n5 1.35656
R1687 ring_out.n7 ring_out.n6 1.35656
R1688 ring_out.n8 ring_out.n7 1.35656
R1689 ring_out.n9 ring_out.n8 1.35656
R1690 ring_out.n10 ring_out.n9 1.35656
R1691 ring_out.n11 ring_out.n10 1.35656
R1692 ring_out.n12 ring_out.n11 1.35656
R1693 ring_out.n13 ring_out.n12 1.35656
R1694 ring_out.n14 ring_out.n13 1.35656
R1695 ring_out.n15 ring_out.n14 0.685584
R1696 ring_out.n2 ring_out.n1 0.303132
R1697 ring_out.n18 ring_out.n2 0.221405
R1698 ring_out.n16 ring_out.n15 0.15724
R1699 ring_out.n18 ring_out.n17 0.0490893
R1700 ring_out ring_out.n18 0.0463464
R1701 ring_out.n17 ring_out.n16 0.0118636
R1702 a_n169_16287.n0 a_n169_16287.n6 113.371
R1703 a_n169_16287.n5 a_n169_16287.n4 113.371
R1704 a_n169_16287.n7 a_n169_16287.t9 74.6407
R1705 a_n169_16287.n2 a_n169_16287.t8 74.6407
R1706 a_n169_16287.t1 a_n169_16287.n3 73.5102
R1707 a_n169_16287.t3 a_n169_16287.n8 73.5102
R1708 a_n169_16287.n4 a_n169_16287.t6 73.5085
R1709 a_n169_16287.n0 a_n169_16287.t3 73.5085
R1710 a_n169_16287.n6 a_n169_16287.t7 73.5085
R1711 a_n169_16287.n5 a_n169_16287.t1 73.5085
R1712 a_n169_16287.n1 a_n169_16287.t0 14.0533
R1713 a_n169_16287.n1 a_n169_16287.t5 11.7371
R1714 a_n169_16287.t4 a_n169_16287.n0 7.79415
R1715 a_n169_16287.n0 a_n169_16287.t2 7.49661
R1716 a_n169_16287.n0 a_n169_16287.n1 5.59997
R1717 a_n169_16287.n8 a_n169_16287.n7 1.13093
R1718 a_n169_16287.n3 a_n169_16287.n2 1.13093
R1719 a_n169_16287.n0 a_n169_16287.n5 0.985754
R1720 a_9754_15288.n0 a_9754_15288.t1 260.2
R1721 a_9754_15288.n1 a_9754_15288.t0 252.136
R1722 a_9754_15288.t4 a_9754_15288.n4 251.333
R1723 a_9754_15288.n2 a_9754_15288.n1 164.748
R1724 a_9754_15288.n4 a_9754_15288.t5 157.893
R1725 a_9754_15288.n3 a_9754_15288.t2 155.667
R1726 a_9754_15288.n0 a_9754_15288.t3 149.827
R1727 a_9754_15288.n3 a_9754_15288.n2 72.9605
R1728 a_9754_15288.n2 a_9754_15288.n0 9.14336
R1729 a_9754_15288.n4 a_9754_15288.n3 8.74717
R1730 a_9754_15288.n1 a_9754_15288.t6 3.16453
R1731 a_5930_14177.n1 a_5930_14177.t1 260.2
R1732 a_5930_14177.n0 a_5930_14177.t0 252.136
R1733 a_5930_14177.t4 a_5930_14177.n4 251.333
R1734 a_5930_14177.n2 a_5930_14177.n0 164.748
R1735 a_5930_14177.n4 a_5930_14177.t6 157.893
R1736 a_5930_14177.n3 a_5930_14177.t2 155.667
R1737 a_5930_14177.n1 a_5930_14177.t3 149.827
R1738 a_5930_14177.n3 a_5930_14177.n2 72.9605
R1739 a_5930_14177.n2 a_5930_14177.n1 9.14336
R1740 a_5930_14177.n4 a_5930_14177.n3 8.74717
R1741 a_5930_14177.n0 a_5930_14177.t5 3.16453
R1742 a_5930_10845.n1 a_5930_10845.t2 260.2
R1743 a_5930_10845.n0 a_5930_10845.t6 252.136
R1744 a_5930_10845.n4 a_5930_10845.t5 251.333
R1745 a_5930_10845.n2 a_5930_10845.n0 164.748
R1746 a_5930_10845.t4 a_5930_10845.n4 157.893
R1747 a_5930_10845.n3 a_5930_10845.t0 155.667
R1748 a_5930_10845.n1 a_5930_10845.t1 149.827
R1749 a_5930_10845.n3 a_5930_10845.n2 72.9605
R1750 a_5930_10845.n2 a_5930_10845.n1 9.14336
R1751 a_5930_10845.n4 a_5930_10845.n3 8.74717
R1752 a_5930_10845.n0 a_5930_10845.t3 3.16453
R1753 ring_100mV_0.mdls_inv_4.IN.n19 ring_100mV_0.mdls_inv_4.IN.t2 265.382
R1754 ring_100mV_0.mdls_inv_4.IN.n21 ring_100mV_0.mdls_inv_4.IN.n20 262.217
R1755 ring_100mV_0.mdls_inv_4.IN.n6 ring_100mV_0.mdls_inv_4.IN.t14 183.099
R1756 ring_100mV_0.mdls_inv_4.IN.n5 ring_100mV_0.mdls_inv_4.IN.t6 183.099
R1757 ring_100mV_0.mdls_inv_4.IN.t6 ring_100mV_0.mdls_inv_4.IN.n4 183.099
R1758 ring_100mV_0.mdls_inv_4.IN.n0 ring_100mV_0.mdls_inv_4.IN.t8 182.653
R1759 ring_100mV_0.mdls_inv_4.IN.t14 ring_100mV_0.mdls_inv_4.IN.n3 182.297
R1760 ring_100mV_0.mdls_inv_4.IN.n0 ring_100mV_0.mdls_inv_4.IN.t11 182.288
R1761 ring_100mV_0.mdls_inv_4.IN.n7 ring_100mV_0.mdls_inv_4.IN.t13 182.285
R1762 ring_100mV_0.mdls_inv_4.IN.n5 ring_100mV_0.mdls_inv_4.IN.t7 182.263
R1763 ring_100mV_0.mdls_inv_4.IN.t13 ring_100mV_0.mdls_inv_4.IN.n6 182.263
R1764 ring_100mV_0.mdls_inv_4.IN.t7 ring_100mV_0.mdls_inv_4.IN.n4 182.263
R1765 ring_100mV_0.mdls_inv_4.IN.n20 ring_100mV_0.mdls_inv_4.IN.t1 155.667
R1766 ring_100mV_0.mdls_inv_4.IN.n19 ring_100mV_0.mdls_inv_4.IN.t0 155.667
R1767 ring_100mV_0.mdls_inv_4.IN.t12 ring_100mV_0.mdls_inv_4.IN.n2 146.282
R1768 ring_100mV_0.mdls_inv_4.IN.n12 ring_100mV_0.mdls_inv_4.IN.t15 145.889
R1769 ring_100mV_0.mdls_inv_4.IN.t15 ring_100mV_0.mdls_inv_4.IN.n11 145.857
R1770 ring_100mV_0.mdls_inv_4.IN.n9 ring_100mV_0.mdls_inv_4.IN.t12 145.851
R1771 ring_100mV_0.mdls_inv_4.IN.n14 ring_100mV_0.mdls_inv_4.IN.t9 135.911
R1772 ring_100mV_0.mdls_inv_4.IN.n17 ring_100mV_0.mdls_inv_4.IN.n16 122.928
R1773 ring_100mV_0.mdls_inv_4.IN.n20 ring_100mV_0.mdls_inv_4.IN.n19 109.715
R1774 ring_100mV_0.mdls_inv_4.IN.t10 ring_100mV_0.mdls_inv_4.IN.n15 98.2234
R1775 ring_100mV_0.mdls_inv_4.IN.n17 ring_100mV_0.mdls_inv_4.IN.t10 49.4098
R1776 ring_100mV_0.mdls_inv_4.IN.n1 ring_100mV_0.mdls_inv_4.IN.t5 45.8204
R1777 ring_100mV_0.mdls_inv_4.IN.n14 ring_100mV_0.mdls_inv_4.IN.n1 28.5785
R1778 ring_100mV_0.mdls_inv_4.IN.n16 ring_100mV_0.mdls_inv_4.IN.t4 28.5685
R1779 ring_100mV_0.mdls_inv_4.IN.t9 ring_100mV_0.mdls_inv_4.IN.n13 19.7637
R1780 ring_100mV_0.mdls_inv_4.IN.n18 ring_100mV_0.mdls_inv_4.IN.n17 5.00095
R1781 ring_100mV_0.mdls_inv_4.IN.n10 ring_100mV_0.mdls_inv_4.IN.n2 4.13208
R1782 ring_100mV_0.mdls_inv_4.IN.n21 ring_100mV_0.mdls_inv_4.IN.t3 3.16453
R1783 ring_100mV_0.mdls_inv_4.IN.n15 ring_100mV_0.mdls_inv_4.IN.n14 2.83669
R1784 ring_100mV_0.mdls_inv_4.IN.n18 ring_100mV_0.mdls_inv_4.IN.n0 1.3453
R1785 ring_100mV_0.mdls_inv_6.OUT ring_100mV_0.mdls_inv_4.IN.n21 1.29092
R1786 ring_100mV_0.mdls_inv_4.IN.n6 ring_100mV_0.mdls_inv_4.IN.n5 0.835457
R1787 ring_100mV_0.mdls_inv_4.IN.n8 ring_100mV_0.mdls_inv_4.IN.n4 0.813812
R1788 ring_100mV_0.mdls_inv_4.IN.n7 ring_100mV_0.mdls_inv_4.IN.n3 0.810242
R1789 ring_100mV_0.mdls_inv_4.IN.n11 ring_100mV_0.mdls_inv_4.IN.n10 0.607643
R1790 ring_100mV_0.mdls_inv_4.IN.n10 ring_100mV_0.mdls_inv_4.IN.n9 0.43198
R1791 ring_100mV_0.mdls_inv_4.IN.n13 ring_100mV_0.mdls_inv_4.IN 0.339159
R1792 ring_100mV_0.mdls_inv_4.IN.n12 ring_100mV_0.mdls_inv_4.IN.n2 0.333833
R1793 ring_100mV_0.mdls_inv_4.IN.n9 ring_100mV_0.mdls_inv_4.IN.n8 0.21421
R1794 ring_100mV_0.mdls_inv_4.IN.n11 ring_100mV_0.mdls_inv_4.IN.n3 0.21421
R1795 ring_100mV_0.mdls_inv_6.OUT ring_100mV_0.mdls_inv_4.IN.n18 0.184521
R1796 ring_100mV_0.mdls_inv_4.IN ring_100mV_0.mdls_inv_4.IN.n12 0.120801
R1797 ring_100mV_0.mdls_inv_4.IN.n8 ring_100mV_0.mdls_inv_4.IN.n7 0.106457
R1798 ldo_out.n9 ldo_out.n8 261.185
R1799 ldo_out.n4 ldo_out.n3 229.173
R1800 ldo_out.n12 ldo_out.n11 74.0415
R1801 ldo_out.n12 ldo_out.n6 72.1843
R1802 ldo_out.n1 ldo_out.t2 7.2144
R1803 ldo_out.n25 ldo_out.t4 5.76538
R1804 ldo_out.n0 ldo_out.t1 4.7068
R1805 ldo_out.n19 ldo_out.t0 4.24157
R1806 ldo_out.n13 ldo_out.n12 1.23559
R1807 ldo_out ldo_out.n25 0.180469
R1808 ldo_out.n24 ldo_out.n23 0.136226
R1809 ldo_out.n24 ldo_out.t3 0.126657
R1810 ldo_out.n14 ldo_out.n1 0.0503555
R1811 ldo_out.n23 ldo_out.n14 0.0427877
R1812 ldo_out.n1 ldo_out.n0 0.0245405
R1813 ldo_out.n25 ldo_out.n24 0.0179077
R1814 ldo_out.n6 ldo_out.n5 0.0153511
R1815 ldo_out.n5 ldo_out.n4 0.014836
R1816 ldo_out.n11 ldo_out.n10 0.0131168
R1817 ldo_out.n10 ldo_out.n9 0.012684
R1818 ldo_out.n21 ldo_out.n20 0.0069195
R1819 ldo_out.n20 ldo_out.n19 0.00641981
R1820 ldo_out.n23 ldo_out.n22 0.00626716
R1821 ldo_out.n21 ldo_out.n16 0.00449474
R1822 ldo_out.n8 ldo_out.n7 0.00432563
R1823 ldo_out.n3 ldo_out.n2 0.00432563
R1824 ldo_out.n16 ldo_out.n15 0.00399493
R1825 ldo_out.n18 ldo_out.n17 0.00345991
R1826 ldo_out.n19 ldo_out.n18 0.00345991
R1827 ldo_out.n22 ldo_out.n21 0.00100012
R1828 ldo_out.n14 ldo_out.n13 0.000504061
R1829 a_n81_16487.t8 a_n81_16487.n4 151.024
R1830 a_n81_16487.t11 a_n81_16487.t7 75.728
R1831 a_n81_16487.t12 a_n81_16487.t8 75.728
R1832 a_n81_16487.t19 a_n81_16487.t12 75.728
R1833 a_n81_16487.t23 a_n81_16487.t19 75.728
R1834 a_n81_16487.t13 a_n81_16487.t23 75.728
R1835 a_n81_16487.t16 a_n81_16487.t13 75.728
R1836 a_n81_16487.t20 a_n81_16487.t16 75.728
R1837 a_n81_16487.t9 a_n81_16487.t20 75.728
R1838 a_n81_16487.t14 a_n81_16487.t9 75.728
R1839 a_n81_16487.t21 a_n81_16487.t14 75.728
R1840 a_n81_16487.t10 a_n81_16487.t21 75.728
R1841 a_n81_16487.t15 a_n81_16487.t10 75.728
R1842 a_n81_16487.t22 a_n81_16487.t15 75.728
R1843 a_n81_16487.t6 a_n81_16487.t22 75.728
R1844 a_n81_16487.t7 a_n81_16487.t17 73.0385
R1845 a_n81_16487.n4 a_n81_16487.t11 61.9359
R1846 a_n81_16487.n1 a_n81_16487.t6 41.3671
R1847 a_n81_16487.n1 a_n81_16487.t0 38.4888
R1848 a_n81_16487.n0 a_n81_16487.t2 37.8394
R1849 a_n81_16487.n5 a_n81_16487.t4 13.5808
R1850 a_n81_16487.n3 a_n81_16487.t1 11.428
R1851 a_n81_16487.n2 a_n81_16487.t3 11.428
R1852 a_n81_16487.n4 a_n81_16487.t18 11.0702
R1853 a_n81_16487.t5 a_n81_16487.n5 10.6813
R1854 a_n81_16487.n5 a_n81_16487.n1 7.30437
R1855 a_n81_16487.n1 a_n81_16487.n3 0.573403
R1856 a_n81_16487.n0 a_n81_16487.n2 0.555619
R1857 a_n81_16487.n3 a_n81_16487.n0 0.403391
R1858 a_3482_8138.n9 a_3482_8138.t15 11.554
R1859 a_3482_8138.n2 a_3482_8138.t14 11.554
R1860 a_3482_8138.n3 a_3482_8138.t12 11.554
R1861 a_3482_8138.n4 a_3482_8138.t19 11.554
R1862 a_3482_8138.n5 a_3482_8138.t16 11.554
R1863 a_3482_8138.n0 a_3482_8138.t10 11.554
R1864 a_3482_8138.n1 a_3482_8138.t17 11.554
R1865 a_3482_8138.n6 a_3482_8138.t13 11.554
R1866 a_3482_8138.n7 a_3482_8138.t11 11.554
R1867 a_3482_8138.n8 a_3482_8138.t18 11.554
R1868 a_3482_8138.n2 a_3482_8138.t8 11.5402
R1869 a_3482_8138.n3 a_3482_8138.t6 11.5402
R1870 a_3482_8138.n4 a_3482_8138.t3 11.5402
R1871 a_3482_8138.n5 a_3482_8138.t0 11.5402
R1872 a_3482_8138.n0 a_3482_8138.t5 11.5402
R1873 a_3482_8138.n1 a_3482_8138.t2 11.5402
R1874 a_3482_8138.n6 a_3482_8138.t7 11.5402
R1875 a_3482_8138.n7 a_3482_8138.t4 11.5402
R1876 a_3482_8138.n8 a_3482_8138.t1 11.5402
R1877 a_3482_8138.t9 a_3482_8138.n9 11.5402
R1878 a_3482_8138.n1 a_3482_8138.n0 7.86782
R1879 a_3482_8138.n3 a_3482_8138.n2 1.26396
R1880 a_3482_8138.n4 a_3482_8138.n3 1.26396
R1881 a_3482_8138.n5 a_3482_8138.n4 1.26396
R1882 a_3482_8138.n7 a_3482_8138.n6 1.26396
R1883 a_3482_8138.n8 a_3482_8138.n7 1.26396
R1884 a_3482_8138.n9 a_3482_8138.n8 1.26396
R1885 a_3482_8138.n6 a_3482_8138.n1 1.26396
R1886 a_3482_8138.n0 a_3482_8138.n5 1.26396
R1887 a_9754_10290.n0 a_9754_10290.t4 260.2
R1888 a_9754_10290.n1 a_9754_10290.t6 252.136
R1889 a_9754_10290.t5 a_9754_10290.n4 251.333
R1890 a_9754_10290.n2 a_9754_10290.n1 164.748
R1891 a_9754_10290.n4 a_9754_10290.t0 157.893
R1892 a_9754_10290.n3 a_9754_10290.t2 155.667
R1893 a_9754_10290.n0 a_9754_10290.t3 149.827
R1894 a_9754_10290.n3 a_9754_10290.n2 72.9605
R1895 a_9754_10290.n2 a_9754_10290.n0 9.14336
R1896 a_9754_10290.n4 a_9754_10290.n3 8.74717
R1897 a_9754_10290.n1 a_9754_10290.t1 3.16453
R1898 a_5930_9179.n1 a_5930_9179.t1 260.2
R1899 a_5930_9179.n0 a_5930_9179.t0 252.136
R1900 a_5930_9179.t4 a_5930_9179.n4 251.333
R1901 a_5930_9179.n2 a_5930_9179.n0 164.748
R1902 a_5930_9179.n4 a_5930_9179.t5 157.893
R1903 a_5930_9179.n3 a_5930_9179.t3 155.667
R1904 a_5930_9179.n1 a_5930_9179.t2 149.827
R1905 a_5930_9179.n3 a_5930_9179.n2 72.9605
R1906 a_5930_9179.n2 a_5930_9179.n1 9.14336
R1907 a_5930_9179.n4 a_5930_9179.n3 8.74717
R1908 a_5930_9179.n0 a_5930_9179.t6 3.16453
R1909 a_5930_12511.t5 a_5930_12511.n4 260.2
R1910 a_5930_12511.n2 a_5930_12511.t6 252.136
R1911 a_5930_12511.n0 a_5930_12511.t2 251.333
R1912 a_5930_12511.n3 a_5930_12511.n2 164.748
R1913 a_5930_12511.n0 a_5930_12511.t0 157.893
R1914 a_5930_12511.n1 a_5930_12511.t3 155.667
R1915 a_5930_12511.n4 a_5930_12511.t4 149.827
R1916 a_5930_12511.n3 a_5930_12511.n1 72.9605
R1917 a_5930_12511.n4 a_5930_12511.n3 9.14336
R1918 a_5930_12511.n1 a_5930_12511.n0 8.74717
R1919 a_5930_12511.n2 a_5930_12511.t1 3.16453
R1920 iref.n0 iref.t1 11.7578
R1921 iref.n0 iref.t0 11.7552
R1922 iref.n1 iref 1.45168
R1923 iref iref.n0 0.151738
R1924 iref.n1 iref 0.0455599
R1925 iref_2nA_0.IREF iref.n1 0.00219179
R1926 ldo_vb.n0 ldo_vb.t1 49.9518
R1927 ldo_vb.n0 ldo_vb.t0 48.1905
R1928 ldo_vb ldo_vb.n0 2.75644
R1929 ldo_vs.n0 ldo_vs.t0 147.147
R1930 ldo_vs.n0 ldo_vs.t1 63.6678
R1931 ldo_vs ldo_vs.n0 44.5008
C0 ring_100mV_0.mdls_inv_2.IN ring_100mV_0.mdls_inv_5.OUT 0.211f
C1 a_9754_7988# ring_100mV_0.mdls_inv_0.OUT 1.21f
C2 ring_100mV_0.mdls_inv_0.IN ring_100mV_0.mdls_inv_0.OUT 2.35f
C3 a_7406_11663# a_9754_11320# 0.0129f
C4 iref_2nA_0.iref_2nA_igenerator_0.Ip2 ring_100mV_0.mdls_inv_1.OUT 3.73e-20
C5 a_1786_16746# iref_2nA_0.iref_2nA_igenerator_0.Vg 0.156f
C6 ldo_vs ldo_iref 0.00227f
C7 a_7406_14995# ring_100mV_0.mdls_inv_2.IN 0.664f
C8 dd_02 a_9754_7988# 1.59f
C9 dd_01 ring_100mV_0.mdls_inv_2.IN 0.0591f
C10 dd_02 ring_100mV_0.mdls_inv_0.IN 4.59f
C11 ring_100mV_0.mdls_inv_1.OUT ring_100mV_0.mdls_inv_7.OUT 0.179f
C12 dd_01 ldo_out 1.37f
C13 a_9754_9654# ring_100mV_0.mdls_inv_1.OUT 0.00146f
C14 ring_100mV_0.mdls_inv_7.OUT ring_100mV_0.mdls_inv_5.OUT 2.1f
C15 a_9754_9654# ring_100mV_0.mdls_inv_5.OUT 1.06e-19
C16 ring_100mV_0.mdls_inv_3.OUT ring_100mV_0.mdls_inv_2.IN 1.46f
C17 a_828_14113# iref 0.143f
C18 iref_2nA_0.iref_2nA_igenerator_0.VCTAT iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.0712f
C19 dd_01 iref_2nA_0.iref_2nA_igenerator_0.Ip2 13.8f
C20 ring_100mV_0.mdls_inv_0.IN ldo_vb 4.67e-20
C21 dd_02 a_9754_11320# 1.59f
C22 ring_100mV_0.mdls_inv_4.IN ring_100mV_0.mdls_inv_5.OUT 0.0308f
C23 ring_100mV_0.mdls_inv_3.OUT iref_2nA_0.iref_2nA_igenerator_0.Ip2 7.84e-20
C24 a_7406_13329# a_9754_12986# 0.0129f
C25 dd_01 ring_100mV_0.mdls_inv_7.OUT 0.144f
C26 dd_02 a_7406_13329# 1.59f
C27 ring_100mV_0.mdls_inv_3.OUT ring_out 0.0153f
C28 iref_2nA_0.iref_2nA_igenerator_0.Ip2 w_583_11504# 0.118f
C29 ring_100mV_0.mdls_inv_0.IN a_9754_7988# 0.669f
C30 ldo_iref ldo_vb 0.267f
C31 ring_100mV_0.mdls_inv_0.OUT a_7406_9997# 2.93e-21
C32 ring_100mV_0.mdls_inv_4.IN a_7406_14995# 1.37e-19
C33 dd_01 ring_100mV_0.mdls_inv_4.IN 0.0221f
C34 ring_100mV_0.mdls_inv_1.OUT ring_100mV_0.mdls_inv_6.IN 1.47f
C35 ring_100mV_0.mdls_inv_2.OUT ring_100mV_0.mdls_inv_5.OUT 2.12f
C36 ring_100mV_0.mdls_inv_5.OUT ring_100mV_0.mdls_inv_6.IN 0.191f
C37 iref_2nA_0.iref_2nA_igenerator_0.Ip2 a_3482_12842# 0.21f
C38 iref_2nA_0.iref_2nA_igenerator_0.Vg iref_2nA_0.iref_2nA_igenerator_0.Ip1 1.14f
C39 iref_2nA_0.iref_2nA_igenerator_0.Ip2 a_3482_12058# 0.361f
C40 ring_100mV_0.mdls_inv_0.IN a_9754_11320# 6.99e-19
C41 dd_02 a_7406_9997# 1.59f
C42 a_9754_14652# ring_100mV_0.mdls_inv_2.IN 0.603f
C43 a_1786_16746# iref_2nA_0.iref_2nA_igenerator_0.Ip1 0.205f
C44 a_1786_15962# dd_01 0.784f
C45 ldo_vs ldo_out 2.36f
C46 ring_100mV_0.mdls_inv_2.OUT a_7406_14995# 6.45e-19
C47 dd_01 ring_100mV_0.mdls_inv_2.OUT 0.132f
C48 dd_01 ring_100mV_0.mdls_inv_6.IN 0.0282f
C49 iref_2nA_0.iref_2nA_igenerator_0.VCTAT iref 0.963f
C50 dd_01 iref 0.815f
C51 a_7406_11663# ring_100mV_0.mdls_inv_7.OUT 6.45e-19
C52 ring_100mV_0.mdls_inv_2.OUT ring_100mV_0.mdls_inv_3.OUT 0.121f
C53 ring_100mV_0.mdls_inv_2.IN a_9754_12986# 1.06e-19
C54 dd_02 ring_100mV_0.mdls_inv_2.IN 6.24f
C55 iref_2nA_0.iref_2nA_igenerator_0.VCTAT a_828_14113# 0.264f
C56 dd_01 a_828_14113# 0.00167f
C57 ring_100mV_0.mdls_inv_0.IN a_7406_9997# 0.00136f
C58 iref w_583_11504# 0.219f
C59 ring_100mV_0.mdls_inv_0.OUT ring_100mV_0.mdls_inv_7.OUT 0.112f
C60 a_9754_9654# ring_100mV_0.mdls_inv_0.OUT 3.31e-19
C61 ring_100mV_0.mdls_inv_4.IN a_7406_11663# 1.07f
C62 ring_100mV_0.mdls_inv_1.OUT a_7406_8331# 1.07f
C63 a_828_14113# w_583_11504# 6.92e-21
C64 iref_2nA_0.iref_2nA_igenerator_0.Vg iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.354f
C65 dd_02 ring_out 1.57f
C66 ldo_vb ldo_out 1.46f
C67 iref a_3482_12842# 0.157f
C68 ring_100mV_0.mdls_inv_7.OUT a_9754_12986# 3.31e-19
C69 dd_02 ring_100mV_0.mdls_inv_7.OUT 4.65f
C70 dd_02 a_9754_9654# 1.59f
C71 a_1786_16746# iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.00404f
C72 a_3482_12058# iref 0.00626f
C73 a_7406_11663# ring_100mV_0.mdls_inv_6.IN 0.664f
C74 dd_01 ring_100mV_0.mdls_inv_1.OUT 0.112f
C75 a_9754_14652# ring_100mV_0.mdls_inv_2.OUT 1.22f
C76 dd_01 ring_100mV_0.mdls_inv_5.OUT 0.144f
C77 ring_100mV_0.mdls_inv_4.IN a_9754_12986# 0.00146f
C78 ring_100mV_0.mdls_inv_4.IN dd_02 4.57f
C79 ldo_vb ring_100mV_0.mdls_inv_7.OUT 0.00182f
C80 ldo_iref ldo_out 0.0248f
C81 a_9754_7988# ring_100mV_0.mdls_inv_7.OUT 1.29e-19
C82 a_7406_13329# ring_100mV_0.mdls_inv_2.IN 1.08f
C83 ring_100mV_0.mdls_inv_0.IN ring_100mV_0.mdls_inv_7.OUT 2.12f
C84 ring_100mV_0.mdls_inv_0.IN a_9754_9654# 1.09f
C85 dd_01 iref_2nA_0.iref_2nA_igenerator_0.VCTAT 0.328f
C86 ring_100mV_0.mdls_inv_2.OUT a_9754_12986# 0.876f
C87 a_1786_15962# iref_2nA_0.iref_2nA_igenerator_0.Vg 0.011f
C88 dd_02 ring_100mV_0.mdls_inv_2.OUT 4.97f
C89 dd_02 ring_100mV_0.mdls_inv_6.IN 4.55f
C90 a_7406_14995# ring_100mV_0.mdls_inv_3.OUT 1.07f
C91 dd_01 ring_100mV_0.mdls_inv_3.OUT 0.00217f
C92 iref_2nA_0.iref_2nA_igenerator_0.VCTAT w_583_11504# 0.228f
C93 iref_2nA_0.iref_2nA_igenerator_0.Vg iref 0.0774f
C94 a_9754_11320# ring_100mV_0.mdls_inv_7.OUT 1.22f
C95 a_1786_15962# a_1786_16746# 1.17f
C96 dd_01 w_583_11504# 1.82f
C97 iref_2nA_0.iref_2nA_igenerator_0.Ip1 iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.493f
C98 iref_2nA_0.iref_2nA_igenerator_0.Vg a_828_14113# 0.785f
C99 a_7406_11663# ring_100mV_0.mdls_inv_1.OUT 1.5e-19
C100 a_7406_11663# ring_100mV_0.mdls_inv_5.OUT 0.00194f
C101 dd_01 vref 1.47f
C102 dd_01 a_3482_12842# 0.51f
C103 a_9754_14652# ring_100mV_0.mdls_inv_5.OUT 0.00215f
C104 ring_100mV_0.mdls_inv_0.IN ring_100mV_0.mdls_inv_6.IN 0.109f
C105 ring_100mV_0.mdls_inv_4.IN a_7406_13329# 0.829f
C106 iref_2nA_0.iref_2nA_igenerator_0.VCTAT a_3482_12058# 3.09e-19
C107 ring_100mV_0.mdls_inv_0.OUT a_7406_8331# 0.607f
C108 dd_01 a_3482_12058# 0.709f
C109 ring_100mV_0.mdls_inv_0.OUT ring_100mV_0.mdls_inv_1.OUT 1.52f
C110 a_7406_9997# ring_100mV_0.mdls_inv_7.OUT 0.00155f
C111 a_9754_9654# a_7406_9997# 0.0129f
C112 a_9754_14652# a_7406_14995# 0.0129f
C113 ring_100mV_0.mdls_inv_2.OUT a_9754_11320# 1.09e-19
C114 a_9754_11320# ring_100mV_0.mdls_inv_6.IN 0.00179f
C115 dd_02 a_7406_8331# 1.59f
C116 dd_02 ring_100mV_0.mdls_inv_1.OUT 4.57f
C117 ring_100mV_0.mdls_inv_5.OUT a_9754_12986# 1.09f
C118 dd_02 ring_100mV_0.mdls_inv_5.OUT 4.62f
C119 ring_100mV_0.mdls_inv_2.IN iref_2nA_0.iref_2nA_igenerator_0.Ip2 9.45e-20
C120 ldo_vs dd_01 0.00151f
C121 ring_100mV_0.mdls_inv_2.OUT a_7406_13329# 0.00155f
C122 a_7406_13329# ring_100mV_0.mdls_inv_6.IN 3.18e-19
C123 dd_01 ring_100mV_0.mdls_inv_0.OUT 0.199f
C124 a_1786_15962# iref_2nA_0.iref_2nA_igenerator_0.Ip1 0.491f
C125 a_3482_12058# a_3482_12842# 1.17f
C126 ldo_vb ring_100mV_0.mdls_inv_5.OUT 6.11e-19
C127 dd_02 a_7406_14995# 1.59f
C128 dd_01 dd_02 0.032f
C129 iref_2nA_0.iref_2nA_igenerator_0.Ip1 iref 0.00398f
C130 a_9754_7988# a_7406_8331# 0.0129f
C131 iref_2nA_0.iref_2nA_igenerator_0.VCTAT iref_2nA_0.iref_2nA_igenerator_0.Vg 0.191f
C132 dd_01 iref_2nA_0.iref_2nA_igenerator_0.Vg 0.511f
C133 ring_100mV_0.mdls_inv_0.IN a_7406_8331# 0.00194f
C134 a_7406_9997# ring_100mV_0.mdls_inv_6.IN 1.07f
C135 ring_100mV_0.mdls_inv_0.IN ring_100mV_0.mdls_inv_1.OUT 0.0308f
C136 ring_100mV_0.mdls_inv_4.IN ring_100mV_0.mdls_inv_2.IN 1.47f
C137 ring_100mV_0.mdls_inv_0.IN ring_100mV_0.mdls_inv_5.OUT 0.134f
C138 dd_02 ring_100mV_0.mdls_inv_3.OUT 4.8f
C139 iref_2nA_0.iref_2nA_igenerator_0.Ip1 a_828_14113# 0.595f
C140 a_1786_16746# dd_01 0.511f
C141 dd_01 ldo_vb 0.0669f
C142 a_9754_9654# ring_100mV_0.mdls_inv_7.OUT 0.876f
C143 ring_100mV_0.mdls_inv_4.IN iref_2nA_0.iref_2nA_igenerator_0.Ip2 1.23e-19
C144 dd_02 vref 0.0607f
C145 a_9754_11320# ring_100mV_0.mdls_inv_5.OUT 0.664f
C146 dd_01 ring_100mV_0.mdls_inv_0.IN 0.172f
C147 ring_100mV_0.mdls_inv_2.OUT ring_100mV_0.mdls_inv_2.IN 1.75f
C148 a_7406_13329# ring_100mV_0.mdls_inv_5.OUT 0.00136f
C149 ring_100mV_0.mdls_inv_4.IN ring_100mV_0.mdls_inv_7.OUT 0.105f
C150 a_1786_15962# iref_2nA_0.iref_2nA_igenerator_0.Ip2 0.00384f
C151 ldo_iref dd_01 0.157f
C152 iref_2nA_0.iref_2nA_igenerator_0.Ip2 ring_100mV_0.mdls_inv_6.IN 1.03e-19
C153 dd_02 a_7406_11663# 1.59f
C154 iref_2nA_0.iref_2nA_igenerator_0.Ip2 iref 1.16f
C155 a_9754_14652# dd_02 1.59f
C156 ring_100mV_0.mdls_inv_1.OUT a_7406_9997# 0.827f
C157 ring_100mV_0.mdls_inv_2.OUT ring_100mV_0.mdls_inv_7.OUT 0.113f
C158 ring_100mV_0.mdls_inv_7.OUT ring_100mV_0.mdls_inv_6.IN 0.015f
C159 iref_2nA_0.iref_2nA_igenerator_0.Ip2 a_828_14113# 0.32f
C160 dd_02 ring_100mV_0.mdls_inv_0.OUT 4.71f
C161 iref_2nA_0.iref_2nA_igenerator_0.VCTAT iref_2nA_0.iref_2nA_igenerator_0.Ip1 0.00286f
C162 dd_01 iref_2nA_0.iref_2nA_igenerator_0.Ip1 6.48f
C163 ring_100mV_0.mdls_inv_4.IN ring_100mV_0.mdls_inv_2.OUT 0.179f
C164 ldo_vs ldo_vb 0.138f
C165 ring_100mV_0.mdls_inv_4.IN ring_100mV_0.mdls_inv_6.IN 1.46f
C166 dd_02 a_9754_12986# 1.59f
C167 ldo_iref ss 9.72f
C168 ldo_vs ss 1.54f
C169 ldo_vb ss 5.33f
C170 vref ss 2.92f
C171 a_9754_7988# ss 0.41f
C172 a_7406_8331# ss 0.41f
C173 ring_100mV_0.mdls_inv_0.OUT ss 8.24f
C174 a_9754_9654# ss 0.41f
C175 ring_100mV_0.mdls_inv_0.IN ss 8.18f
C176 a_7406_9997# ss 0.41f
C177 ring_100mV_0.mdls_inv_1.OUT ss 8.17f
C178 a_9754_11320# ss 0.41f
C179 ring_100mV_0.mdls_inv_7.OUT ss 8.13f
C180 a_7406_11663# ss 0.41f
C181 ring_100mV_0.mdls_inv_6.IN ss 8.5f
C182 a_9754_12986# ss 0.41f
C183 ring_100mV_0.mdls_inv_5.OUT ss 8.14f
C184 a_7406_13329# ss 0.41f
C185 ring_100mV_0.mdls_inv_4.IN ss 8.22f
C186 a_9754_14652# ss 0.41f
C187 ring_100mV_0.mdls_inv_2.OUT ss 8.09f
C188 a_7406_14995# ss 0.41f
C189 ring_100mV_0.mdls_inv_2.IN ss 13f
C190 ring_100mV_0.mdls_inv_3.OUT ss 13f
C191 ring_out ss 22.5f
C192 a_3482_12842# ss 0.267f
C193 iref ss 6.88f
C194 a_3482_12058# ss 0.339f
C195 a_828_14113# ss 0.955f
C196 iref_2nA_0.iref_2nA_igenerator_0.Ip2 ss 9.88f
C197 a_1786_16746# ss 0.267f
C198 a_1786_15962# ss 0.31f
C199 iref_2nA_0.iref_2nA_igenerator_0.Ip1 ss 3.65f
C200 iref_2nA_0.iref_2nA_igenerator_0.Vg ss 7.52f
C201 ldo_out ss 12f
C202 w_583_11504# ss 6.69f
C203 iref_2nA_0.iref_2nA_igenerator_0.VCTAT ss 13.6f
C204 dd_02 ss 71.9f
C205 dd_01 ss 0.176p
C206 ldo_vs.t1 ss 0.764f
C207 ldo_vs.t0 ss 0.947f
C208 ldo_vs.n0 ss 6.9e-19
C209 ldo_vb.t0 ss 0.246f
C210 ldo_vb.t1 ss 0.263f
C211 ldo_vb.n0 ss 1.68f
C212 iref.t0 ss 0.0062f
C213 iref.t1 ss 0.00622f
C214 iref.n0 ss 0.159f
C215 iref.n1 ss 1.15f
C216 iref_2nA_0.IREF ss 0.415f
C217 a_5930_12511.t3 ss 0.95f
C218 a_5930_12511.t0 ss 0.939f
C219 a_5930_12511.t2 ss 1.01f
C220 a_5930_12511.n0 ss 0.244f
C221 a_5930_12511.n1 ss 0.172f
C222 a_5930_12511.t6 ss 0.451f
C223 a_5930_12511.t1 ss 0.0858f
C224 a_5930_12511.n2 ss 0.91f
C225 a_5930_12511.n3 ss 0.154f
C226 a_5930_12511.t4 ss 0.946f
C227 a_5930_12511.n4 ss 0.234f
C228 a_5930_12511.t5 ss 1.01f
C229 a_5930_9179.t5 ss 0.939f
C230 a_5930_9179.t3 ss 0.95f
C231 a_5930_9179.t0 ss 0.451f
C232 a_5930_9179.t6 ss 0.0858f
C233 a_5930_9179.n0 ss 0.91f
C234 a_5930_9179.t1 ss 1.01f
C235 a_5930_9179.t2 ss 0.946f
C236 a_5930_9179.n1 ss 0.234f
C237 a_5930_9179.n2 ss 0.154f
C238 a_5930_9179.n3 ss 0.172f
C239 a_5930_9179.n4 ss 0.244f
C240 a_5930_9179.t4 ss 1.01f
C241 a_9754_10290.t0 ss 0.939f
C242 a_9754_10290.t2 ss 0.95f
C243 a_9754_10290.t4 ss 1.01f
C244 a_9754_10290.t3 ss 0.946f
C245 a_9754_10290.n0 ss 0.234f
C246 a_9754_10290.t6 ss 0.451f
C247 a_9754_10290.t1 ss 0.0858f
C248 a_9754_10290.n1 ss 0.91f
C249 a_9754_10290.n2 ss 0.154f
C250 a_9754_10290.n3 ss 0.172f
C251 a_9754_10290.n4 ss 0.244f
C252 a_9754_10290.t5 ss 1.01f
C253 a_3482_8138.n0 ss 0.9f
C254 a_3482_8138.n1 ss 0.9f
C255 a_3482_8138.t17 ss 0.028f
C256 a_3482_8138.t2 ss 0.0279f
C257 a_3482_8138.t14 ss 0.028f
C258 a_3482_8138.t8 ss 0.0279f
C259 a_3482_8138.n2 ss 0.372f
C260 a_3482_8138.t12 ss 0.028f
C261 a_3482_8138.t6 ss 0.0279f
C262 a_3482_8138.n3 ss 0.45f
C263 a_3482_8138.t19 ss 0.028f
C264 a_3482_8138.t3 ss 0.0279f
C265 a_3482_8138.n4 ss 0.45f
C266 a_3482_8138.t16 ss 0.028f
C267 a_3482_8138.t0 ss 0.0279f
C268 a_3482_8138.n5 ss 0.448f
C269 a_3482_8138.t10 ss 0.028f
C270 a_3482_8138.t5 ss 0.0279f
C271 a_3482_8138.t13 ss 0.028f
C272 a_3482_8138.t7 ss 0.0279f
C273 a_3482_8138.n6 ss 0.448f
C274 a_3482_8138.t11 ss 0.028f
C275 a_3482_8138.t4 ss 0.0279f
C276 a_3482_8138.n7 ss 0.45f
C277 a_3482_8138.t18 ss 0.028f
C278 a_3482_8138.t1 ss 0.0279f
C279 a_3482_8138.n8 ss 0.45f
C280 a_3482_8138.t15 ss 0.028f
C281 a_3482_8138.n9 ss 0.372f
C282 a_3482_8138.t9 ss 0.0279f
C283 a_n81_16487.n0 ss 0.731f
C284 a_n81_16487.n1 ss 3.4f
C285 a_n81_16487.t0 ss 0.305f
C286 a_n81_16487.t3 ss 0.0174f
C287 a_n81_16487.n2 ss 0.447f
C288 a_n81_16487.t2 ss 0.309f
C289 a_n81_16487.t1 ss 0.0174f
C290 a_n81_16487.n3 ss 0.156f
C291 a_n81_16487.t17 ss 0.92f
C292 a_n81_16487.t7 ss 0.935f
C293 a_n81_16487.t11 ss 0.858f
C294 a_n81_16487.t18 ss 0.492f
C295 a_n81_16487.n4 ss 0.828f
C296 a_n81_16487.t8 ss 1.68f
C297 a_n81_16487.t12 ss 0.919f
C298 a_n81_16487.t19 ss 0.919f
C299 a_n81_16487.t23 ss 0.919f
C300 a_n81_16487.t13 ss 0.919f
C301 a_n81_16487.t16 ss 0.919f
C302 a_n81_16487.t20 ss 0.919f
C303 a_n81_16487.t9 ss 0.919f
C304 a_n81_16487.t14 ss 0.919f
C305 a_n81_16487.t21 ss 0.919f
C306 a_n81_16487.t10 ss 0.919f
C307 a_n81_16487.t15 ss 0.919f
C308 a_n81_16487.t22 ss 0.919f
C309 a_n81_16487.t6 ss 0.65f
C310 a_n81_16487.t4 ss 0.226f
C311 a_n81_16487.n5 ss 2.78f
C312 a_n81_16487.t5 ss 0.13f
C313 ldo_out.t4 ss 0.0258f
C314 ldo_out.t3 ss 4.98f
C315 ldo_out.t2 ss 0.161f
C316 ldo_out.t1 ss 0.0261f
C317 ldo_out.n0 ss 0.108f
C318 ldo_out.n1 ss 0.408f
C319 ldo_out.n2 ss 0.0596f
C320 ldo_out.n3 ss 0.512f
C321 ldo_out.n4 ss 0.728f
C322 ldo_out.n5 ss 0.0341f
C323 ldo_out.n6 ss 0.0305f
C324 ldo_out.n7 ss 0.061f
C325 ldo_out.n8 ss 0.564f
C326 ldo_out.n9 ss 0.78f
C327 ldo_out.n10 ss 0.0354f
C328 ldo_out.n11 ss 0.0318f
C329 ldo_out.n12 ss 0.0562f
C330 ldo_out.n13 ss 0.0137f
C331 ldo_out.n14 ss 0.00788f
C332 ldo_out.n15 ss 0.426f
C333 ldo_out.n16 ss 0.0109f
C334 ldo_out.n17 ss 0.0705f
C335 ldo_out.n18 ss 0.0705f
C336 ldo_out.t0 ss 0.0508f
C337 ldo_out.n19 ss 0.388f
C338 ldo_out.n20 ss 0.011f
C339 ldo_out.n22 ss 0.0367f
C340 ldo_out.n23 ss 0.0359f
C341 ldo_out.n24 ss 1.44f
C342 ldo_out.n25 ss 0.305f
C343 ring_100mV_0.mdls_inv_4.IN.t8 ss 0.153f
C344 ring_100mV_0.mdls_inv_4.IN.t11 ss 0.152f
C345 ring_100mV_0.mdls_inv_4.IN.n0 ss 0.445f
C346 ring_100mV_0.mdls_inv_4.IN.t5 ss 0.196f
C347 ring_100mV_0.mdls_inv_4.IN.n1 ss 0.0764f
C348 ring_100mV_0.mdls_inv_4.IN.n2 ss 0.377f
C349 ring_100mV_0.mdls_inv_4.IN.n3 ss 0.251f
C350 ring_100mV_0.mdls_inv_4.IN.n4 ss 0.488f
C351 ring_100mV_0.mdls_inv_4.IN.t6 ss 0.302f
C352 ring_100mV_0.mdls_inv_4.IN.t7 ss 0.3f
C353 ring_100mV_0.mdls_inv_4.IN.n5 ss 0.489f
C354 ring_100mV_0.mdls_inv_4.IN.t14 ss 0.301f
C355 ring_100mV_0.mdls_inv_4.IN.n6 ss 0.489f
C356 ring_100mV_0.mdls_inv_4.IN.t13 ss 0.3f
C357 ring_100mV_0.mdls_inv_4.IN.n7 ss 0.227f
C358 ring_100mV_0.mdls_inv_4.IN.n8 ss 0.0354f
C359 ring_100mV_0.mdls_inv_4.IN.t12 ss 0.376f
C360 ring_100mV_0.mdls_inv_4.IN.n9 ss 0.296f
C361 ring_100mV_0.mdls_inv_4.IN.n10 ss 0.0983f
C362 ring_100mV_0.mdls_inv_4.IN.n11 ss 0.294f
C363 ring_100mV_0.mdls_inv_4.IN.t15 ss 0.376f
C364 ring_100mV_0.mdls_inv_4.IN.n12 ss 0.307f
C365 ring_100mV_0.mdls_inv_4.IN.n13 ss 0.282f
C366 ring_100mV_0.mdls_inv_4.IN.t9 ss 0.406f
C367 ring_100mV_0.mdls_inv_4.IN.n14 ss 0.64f
C368 ring_100mV_0.mdls_inv_4.IN.n15 ss 0.605f
C369 ring_100mV_0.mdls_inv_4.IN.t10 ss 0.14f
C370 ring_100mV_0.mdls_inv_4.IN.t4 ss 0.009f
C371 ring_100mV_0.mdls_inv_4.IN.n16 ss 0.103f
C372 ring_100mV_0.mdls_inv_4.IN.n17 ss 0.265f
C373 ring_100mV_0.mdls_inv_4.IN.n18 ss 0.376f
C374 ring_100mV_0.mdls_inv_4.IN.t1 ss 0.548f
C375 ring_100mV_0.mdls_inv_4.IN.t0 ss 0.548f
C376 ring_100mV_0.mdls_inv_4.IN.t2 ss 0.585f
C377 ring_100mV_0.mdls_inv_4.IN.n19 ss 0.163f
C378 ring_100mV_0.mdls_inv_4.IN.n20 ss 0.157f
C379 ring_100mV_0.mdls_inv_4.IN.t3 ss 0.0495f
C380 ring_100mV_0.mdls_inv_4.IN.n21 ss 0.412f
C381 ring_100mV_0.mdls_inv_6.OUT ss 0.0825f
C382 a_5930_10845.t0 ss 0.963f
C383 a_5930_10845.t6 ss 0.458f
C384 a_5930_10845.t3 ss 0.087f
C385 a_5930_10845.n0 ss 0.923f
C386 a_5930_10845.t2 ss 1.02f
C387 a_5930_10845.t1 ss 0.959f
C388 a_5930_10845.n1 ss 0.238f
C389 a_5930_10845.n2 ss 0.156f
C390 a_5930_10845.n3 ss 0.175f
C391 a_5930_10845.t5 ss 1.02f
C392 a_5930_10845.n4 ss 0.247f
C393 a_5930_10845.t4 ss 0.952f
C394 a_5930_14177.t6 ss 0.952f
C395 a_5930_14177.t2 ss 0.963f
C396 a_5930_14177.t0 ss 0.458f
C397 a_5930_14177.t5 ss 0.087f
C398 a_5930_14177.n0 ss 0.923f
C399 a_5930_14177.t1 ss 1.02f
C400 a_5930_14177.t3 ss 0.959f
C401 a_5930_14177.n1 ss 0.238f
C402 a_5930_14177.n2 ss 0.156f
C403 a_5930_14177.n3 ss 0.175f
C404 a_5930_14177.n4 ss 0.247f
C405 a_5930_14177.t4 ss 1.02f
C406 a_9754_15288.t5 ss 0.939f
C407 a_9754_15288.t2 ss 0.95f
C408 a_9754_15288.t1 ss 1.01f
C409 a_9754_15288.t3 ss 0.946f
C410 a_9754_15288.n0 ss 0.234f
C411 a_9754_15288.t0 ss 0.451f
C412 a_9754_15288.t6 ss 0.0858f
C413 a_9754_15288.n1 ss 0.91f
C414 a_9754_15288.n2 ss 0.154f
C415 a_9754_15288.n3 ss 0.172f
C416 a_9754_15288.n4 ss 0.244f
C417 a_9754_15288.t4 ss 1.01f
C418 a_n169_16287.n0 ss 0.606f
C419 a_n169_16287.t5 ss 0.00857f
C420 a_n169_16287.t0 ss 0.0398f
C421 a_n169_16287.n1 ss 0.702f
C422 a_n169_16287.t2 ss 0.0133f
C423 a_n169_16287.t8 ss 0.104f
C424 a_n169_16287.n2 ss 0.125f
C425 a_n169_16287.n3 ss 0.0654f
C426 a_n169_16287.t1 ss 0.0633f
C427 a_n169_16287.t6 ss 0.0633f
C428 a_n169_16287.n4 ss 0.0962f
C429 a_n169_16287.n5 ss 0.0792f
C430 a_n169_16287.t7 ss 0.0633f
C431 a_n169_16287.n6 ss 0.0962f
C432 a_n169_16287.t9 ss 0.104f
C433 a_n169_16287.n7 ss 0.125f
C434 a_n169_16287.n8 ss 0.0654f
C435 a_n169_16287.t3 ss 0.0633f
C436 a_n169_16287.t4 ss 0.0168f
C437 ring_out.t9 ss 0.0895f
C438 ring_out.t1 ss 0.0076f
C439 ring_out.t3 ss 0.00508f
C440 ring_out.n0 ss 0.145f
C441 ring_out.t0 ss 0.00508f
C442 ring_out.n1 ss 0.0753f
C443 ring_out.t2 ss 0.00607f
C444 ring_out.n2 ss 0.0841f
C445 ring_out.t19 ss 0.0882f
C446 ring_out.t13 ss 0.0882f
C447 ring_out.t10 ss 0.136f
C448 ring_out.t17 ss 0.0904f
C449 ring_out.n3 ss 0.359f
C450 ring_out.t7 ss 0.0904f
C451 ring_out.n4 ss 0.206f
C452 ring_out.t14 ss 0.0904f
C453 ring_out.n5 ss 0.206f
C454 ring_out.t4 ss 0.0904f
C455 ring_out.n6 ss 0.206f
C456 ring_out.t11 ss 0.0904f
C457 ring_out.n7 ss 0.206f
C458 ring_out.t18 ss 0.0904f
C459 ring_out.n8 ss 0.206f
C460 ring_out.t8 ss 0.0904f
C461 ring_out.n9 ss 0.206f
C462 ring_out.t15 ss 0.0904f
C463 ring_out.n10 ss 0.206f
C464 ring_out.t5 ss 0.0904f
C465 ring_out.n11 ss 0.206f
C466 ring_out.t12 ss 0.0904f
C467 ring_out.n12 ss 0.206f
C468 ring_out.t16 ss 0.0904f
C469 ring_out.n13 ss 0.206f
C470 ring_out.t6 ss 0.0904f
C471 ring_out.n14 ss 0.208f
C472 ring_out.n15 ss 0.37f
C473 ring_out.n16 ss 0.283f
C474 ring_out.n17 ss 0.859f
C475 ring_out.n18 ss 0.0683f
C476 a_5712_16467.t5 ss 0.205f
C477 a_5712_16467.t8 ss 0.139f
C478 a_5712_16467.n0 ss 0.527f
C479 a_5712_16467.t3 ss 0.139f
C480 a_5712_16467.n1 ss 0.303f
C481 a_5712_16467.t7 ss 0.139f
C482 a_5712_16467.n2 ss 0.303f
C483 a_5712_16467.t2 ss 0.139f
C484 a_5712_16467.n3 ss 0.303f
C485 a_5712_16467.t6 ss 0.139f
C486 a_5712_16467.n4 ss 0.303f
C487 a_5712_16467.t21 ss 0.194f
C488 a_5712_16467.n5 ss 0.251f
C489 a_5712_16467.t12 ss 0.194f
C490 a_5712_16467.n6 ss 0.263f
C491 a_5712_16467.t25 ss 0.194f
C492 a_5712_16467.n7 ss 0.149f
C493 a_5712_16467.t16 ss 0.194f
C494 a_5712_16467.n8 ss 0.149f
C495 a_5712_16467.t29 ss 0.194f
C496 a_5712_16467.n9 ss 0.149f
C497 a_5712_16467.t20 ss 0.194f
C498 a_5712_16467.n10 ss 0.149f
C499 a_5712_16467.n11 ss 0.267f
C500 a_5712_16467.n12 ss 0.149f
C501 a_5712_16467.n13 ss 0.149f
C502 a_5712_16467.n14 ss 0.149f
C503 a_5712_16467.n15 ss 0.149f
C504 a_5712_16467.n16 ss 0.149f
C505 a_5712_16467.t11 ss 0.194f
C506 a_5712_16467.n17 ss 0.149f
C507 a_5712_16467.t23 ss 0.194f
C508 a_5712_16467.n18 ss 0.149f
C509 a_5712_16467.n19 ss 0.149f
C510 a_5712_16467.n20 ss 0.149f
C511 a_5712_16467.t14 ss 0.194f
C512 a_5712_16467.n21 ss 0.149f
C513 a_5712_16467.t27 ss 0.194f
C514 a_5712_16467.n22 ss 0.149f
C515 a_5712_16467.n23 ss 0.149f
C516 a_5712_16467.n24 ss 0.149f
C517 a_5712_16467.t18 ss 0.194f
C518 a_5712_16467.n25 ss 0.139f
C519 a_5712_16467.t22 ss 0.322f
C520 a_5712_16467.t10 ss 0.194f
C521 a_5712_16467.n26 ss 0.226f
C522 a_5712_16467.t17 ss 0.194f
C523 a_5712_16467.n27 ss 0.149f
C524 a_5712_16467.t26 ss 0.194f
C525 a_5712_16467.n28 ss 0.149f
C526 a_5712_16467.n29 ss 0.226f
C527 a_5712_16467.n30 ss 0.149f
C528 a_5712_16467.n31 ss 0.149f
C529 a_5712_16467.n32 ss 0.149f
C530 a_5712_16467.t13 ss 0.194f
C531 a_5712_16467.n33 ss 0.14f
C532 a_5712_16467.n34 ss 0.104f
C533 a_5712_16467.t1 ss 0.00583f
C534 a_5712_16467.t19 ss 0.125f
C535 a_5712_16467.n35 ss 0.0749f
C536 a_5712_16467.t28 ss 0.0527f
C537 a_5712_16467.n36 ss 0.0889f
C538 a_5712_16467.t15 ss 0.0527f
C539 a_5712_16467.n37 ss 0.0707f
C540 a_5712_16467.n38 ss 0.0889f
C541 a_5712_16467.n39 ss 0.0707f
C542 a_5712_16467.n40 ss 0.0561f
C543 a_5712_16467.n41 ss 0.0295f
C544 a_5712_16467.t24 ss 0.0885f
C545 a_5712_16467.n42 ss 0.0928f
C546 a_5712_16467.n43 ss 0.139f
C547 a_5712_16467.t0 ss 0.011f
C548 a_5712_16467.n44 ss 0.568f
C549 a_5712_16467.t4 ss 0.139f
C550 a_5712_16467.n45 ss 0.327f
C551 a_5712_16467.n46 ss 0.303f
C552 a_5712_16467.t9 ss 0.139f
C553 a_955_10311.t2 ss 0.845f
C554 a_955_10311.t1 ss 0.0037f
C555 a_955_10311.n0 ss 1.41f
C556 a_955_10311.t0 ss 0.0412f
C557 a_9754_11956.t5 ss 0.939f
C558 a_9754_11956.t2 ss 0.95f
C559 a_9754_11956.t1 ss 1.01f
C560 a_9754_11956.t3 ss 0.946f
C561 a_9754_11956.n0 ss 0.234f
C562 a_9754_11956.t0 ss 0.451f
C563 a_9754_11956.t6 ss 0.0858f
C564 a_9754_11956.n1 ss 0.91f
C565 a_9754_11956.n2 ss 0.154f
C566 a_9754_11956.n3 ss 0.172f
C567 a_9754_11956.n4 ss 0.244f
C568 a_9754_11956.t4 ss 1.01f
C569 a_5930_7513.t6 ss 0.451f
C570 a_5930_7513.t5 ss 0.0858f
C571 a_5930_7513.n0 ss 0.91f
C572 a_5930_7513.t1 ss 1.01f
C573 a_5930_7513.t0 ss 0.946f
C574 a_5930_7513.n1 ss 0.234f
C575 a_5930_7513.n2 ss 0.154f
C576 a_5930_7513.t4 ss 0.939f
C577 a_5930_7513.t2 ss 1.01f
C578 a_5930_7513.n3 ss 0.244f
C579 a_5930_7513.n4 ss 0.172f
C580 a_5930_7513.t3 ss 0.95f
C581 a_14490_9380.n0 ss 0.805f
C582 a_14490_9380.t4 ss 0.0697f
C583 a_14490_9380.t0 ss 0.00837f
C584 a_14490_9380.t1 ss 0.00533f
C585 a_14490_9380.t5 ss 7.79f
C586 a_14490_9380.t3 ss 0.0231f
C587 a_14490_9380.n1 ss 0.898f
C588 a_14490_9380.t2 ss 0.1f
C589 a_15054_7578.n0 ss 0.0881f
C590 a_15054_7578.n1 ss 0.941f
C591 a_15054_7578.t4 ss 0.351f
C592 a_15054_7578.t6 ss 0.719f
C593 a_15054_7578.t0 ss 0.429f
C594 a_15054_7578.n2 ss 0.229f
C595 a_15054_7578.t1 ss 0.00554f
C596 a_15054_7578.t7 ss 0.719f
C597 a_15054_7578.t2 ss 0.429f
C598 a_15054_7578.n3 ss 0.229f
C599 a_15054_7578.t3 ss 0.00554f
C600 a_15054_7578.n4 ss 1.09f
C601 a_15054_7578.t5 ss 0.162f
C602 ring_100mV_0.mdls_inv_8.IN ss 0.407f
C603 ring_100mV_0.mdls_inv_1.OUT.n0 ss 0.251f
C604 ring_100mV_0.mdls_inv_1.OUT.n1 ss 0.263f
C605 ring_100mV_0.mdls_inv_1.OUT.t9 ss 0.153f
C606 ring_100mV_0.mdls_inv_1.OUT.t15 ss 0.152f
C607 ring_100mV_0.mdls_inv_1.OUT.n2 ss 0.445f
C608 ring_100mV_0.mdls_inv_1.OUT.t6 ss 0.196f
C609 ring_100mV_0.mdls_inv_1.OUT.n3 ss 0.0764f
C610 ring_100mV_0.mdls_inv_1.OUT.n4 ss 0.377f
C611 ring_100mV_0.mdls_inv_1.OUT.n5 ss 0.488f
C612 ring_100mV_0.mdls_inv_1.OUT.t11 ss 0.302f
C613 ring_100mV_0.mdls_inv_1.OUT.t8 ss 0.3f
C614 ring_100mV_0.mdls_inv_1.OUT.n6 ss 0.489f
C615 ring_100mV_0.mdls_inv_1.OUT.t5 ss 0.301f
C616 ring_100mV_0.mdls_inv_1.OUT.n7 ss 0.489f
C617 ring_100mV_0.mdls_inv_1.OUT.t7 ss 0.3f
C618 ring_100mV_0.mdls_inv_1.OUT.t10 ss 0.376f
C619 ring_100mV_0.mdls_inv_1.OUT.n8 ss 0.295f
C620 ring_100mV_0.mdls_inv_1.OUT.n9 ss 0.0983f
C621 ring_100mV_0.mdls_inv_1.OUT.n10 ss 0.294f
C622 ring_100mV_0.mdls_inv_1.OUT.t13 ss 0.376f
C623 ring_100mV_0.mdls_inv_1.OUT.n11 ss 0.282f
C624 ring_100mV_0.mdls_inv_1.OUT.t12 ss 0.406f
C625 ring_100mV_0.mdls_inv_1.OUT.n12 ss 0.641f
C626 ring_100mV_0.mdls_inv_1.OUT.n13 ss 0.606f
C627 ring_100mV_0.mdls_inv_1.OUT.t14 ss 0.14f
C628 ring_100mV_0.mdls_inv_1.OUT.t2 ss 0.009f
C629 ring_100mV_0.mdls_inv_1.OUT.n14 ss 0.103f
C630 ring_100mV_0.mdls_inv_1.OUT.n15 ss 0.265f
C631 ring_100mV_0.mdls_inv_1.OUT.n16 ss 0.376f
C632 ring_100mV_0.mdls_inv_1.OUT.t4 ss 0.548f
C633 ring_100mV_0.mdls_inv_1.OUT.t3 ss 0.585f
C634 ring_100mV_0.mdls_inv_1.OUT.n17 ss 0.163f
C635 ring_100mV_0.mdls_inv_1.OUT.t0 ss 0.548f
C636 ring_100mV_0.mdls_inv_1.OUT.n18 ss 0.157f
C637 ring_100mV_0.mdls_inv_1.OUT.t1 ss 0.0495f
C638 ring_100mV_0.mdls_inv_1.OUT.n19 ss 0.412f
C639 ring_100mV_0.mdls_inv_0.OUT.t0 ss 0.652f
C640 ring_100mV_0.mdls_inv_0.OUT.t2 ss 0.696f
C641 ring_100mV_0.mdls_inv_0.OUT.t3 ss 0.652f
C642 ring_100mV_0.mdls_inv_0.OUT.n0 ss 0.194f
C643 ring_100mV_0.mdls_inv_0.OUT.n1 ss 0.186f
C644 ring_100mV_0.mdls_inv_0.OUT.t1 ss 0.0589f
C645 ring_100mV_0.mdls_inv_0.OUT.n2 ss 0.494f
C646 ring_100mV_0.mdls_inv_0.OUT.t9 ss 0.181f
C647 ring_100mV_0.mdls_inv_0.OUT.t15 ss 0.182f
C648 ring_100mV_0.mdls_inv_0.OUT.n3 ss 0.529f
C649 ring_100mV_0.mdls_inv_0.OUT.t5 ss 0.233f
C650 ring_100mV_0.mdls_inv_0.OUT.n4 ss 0.0909f
C651 ring_100mV_0.mdls_inv_0.OUT.n5 ss 0.448f
C652 ring_100mV_0.mdls_inv_0.OUT.n6 ss 0.299f
C653 ring_100mV_0.mdls_inv_0.OUT.n7 ss 0.58f
C654 ring_100mV_0.mdls_inv_0.OUT.t12 ss 0.36f
C655 ring_100mV_0.mdls_inv_0.OUT.t13 ss 0.357f
C656 ring_100mV_0.mdls_inv_0.OUT.n8 ss 0.582f
C657 ring_100mV_0.mdls_inv_0.OUT.t7 ss 0.358f
C658 ring_100mV_0.mdls_inv_0.OUT.n9 ss 0.582f
C659 ring_100mV_0.mdls_inv_0.OUT.t6 ss 0.357f
C660 ring_100mV_0.mdls_inv_0.OUT.n10 ss 0.27f
C661 ring_100mV_0.mdls_inv_0.OUT.n11 ss 0.0421f
C662 ring_100mV_0.mdls_inv_0.OUT.t8 ss 0.448f
C663 ring_100mV_0.mdls_inv_0.OUT.n12 ss 0.351f
C664 ring_100mV_0.mdls_inv_0.OUT.n13 ss 0.117f
C665 ring_100mV_0.mdls_inv_0.OUT.n14 ss 0.35f
C666 ring_100mV_0.mdls_inv_0.OUT.t14 ss 0.447f
C667 ring_100mV_0.mdls_inv_0.OUT.n15 ss 0.366f
C668 ring_100mV_0.mdls_inv_1.IN ss 0.118f
C669 ring_100mV_0.mdls_inv_0.OUT.n16 ss 0.335f
C670 ring_100mV_0.mdls_inv_0.OUT.t11 ss 0.482f
C671 ring_100mV_0.mdls_inv_0.OUT.n17 ss 0.801f
C672 ring_100mV_0.mdls_inv_0.OUT.n18 ss 0.847f
C673 ring_100mV_0.mdls_inv_0.OUT.t10 ss 0.166f
C674 ring_100mV_0.mdls_inv_0.OUT.t4 ss 0.0107f
C675 ring_100mV_0.mdls_inv_0.OUT.n19 ss 0.123f
C676 ring_100mV_0.mdls_inv_0.OUT.n20 ss 0.315f
C677 ring_100mV_0.mdls_inv_0.OUT.n21 ss 0.441f
C678 a_9754_8624.t1 ss 0.95f
C679 a_9754_8624.t3 ss 0.939f
C680 a_9754_8624.t2 ss 1.01f
C681 a_9754_8624.n0 ss 0.244f
C682 a_9754_8624.n1 ss 0.172f
C683 a_9754_8624.t6 ss 1.01f
C684 a_9754_8624.t5 ss 0.946f
C685 a_9754_8624.n2 ss 0.234f
C686 a_9754_8624.n3 ss 0.154f
C687 a_9754_8624.t0 ss 0.451f
C688 a_9754_8624.n4 ss 0.91f
C689 a_9754_8624.t4 ss 0.0858f
C690 a_14834_9380.t2 ss 0.228f
C691 a_14834_9380.t3 ss 0.0347f
C692 a_14834_9380.n0 ss 0.868f
C693 a_14834_9380.t7 ss 0.102f
C694 a_14834_9380.t4 ss 0.102f
C695 a_14834_9380.t1 ss 0.144f
C696 a_14834_9380.t0 ss 0.12f
C697 a_14834_9380.n1 ss 1.39f
C698 a_14834_9380.t5 ss 0.113f
C699 a_14834_9380.n2 ss 0.748f
C700 a_14834_9380.n3 ss 0.386f
C701 a_14834_9380.n4 ss 0.385f
C702 a_14834_9380.n5 ss 0.664f
C703 a_14834_9380.t6 ss 0.114f
C704 a_16150_16902.n0 ss 0.358f
C705 a_16150_16902.t4 ss 0.131f
C706 a_16150_16902.t2 ss 0.13f
C707 a_16150_16902.t6 ss 0.0352f
C708 a_16150_16902.t0 ss 0.157f
C709 a_16150_16902.t3 ss 0.0194f
C710 a_16150_16902.n1 ss 0.251f
C711 a_16150_16902.n2 ss 0.291f
C712 a_16150_16902.t1 ss 0.00621f
C713 a_16150_16902.n3 ss 0.126f
C714 a_16150_16902.n4 ss 0.0485f
C715 a_16150_16902.n5 ss 0.095f
C716 a_16150_16902.n6 ss 0.164f
C717 a_16150_16902.n7 ss 0.305f
C718 a_16150_16902.t5 ss 0.0832f
C719 ring_100mV_0.mdls_inv_3.OUT.n0 ss 1.59f
C720 ring_100mV_0.mdls_inv_3.OUT.t5 ss 0.13f
C721 ring_100mV_0.mdls_inv_3.OUT.t10 ss 0.129f
C722 ring_100mV_0.mdls_inv_3.OUT.n1 ss 0.378f
C723 ring_100mV_0.ring_100mV_buffer_0.IN ss 0.443f
C724 ring_100mV_0.mdls_inv_3.OUT.t6 ss 0.164f
C725 ring_100mV_0.mdls_inv_3.OUT.t11 ss 0.176f
C726 ring_100mV_0.mdls_inv_3.OUT.n2 ss 0.0691f
C727 ring_100mV_0.mdls_inv_3.OUT.n3 ss 0.387f
C728 ring_100mV_0.mdls_inv_3.OUT.n4 ss 0.235f
C729 ring_100mV_0.mdls_inv_3.OUT.n5 ss 0.235f
C730 ring_100mV_0.mdls_inv_3.OUT.n6 ss 0.235f
C731 ring_100mV_0.mdls_inv_3.OUT.n7 ss 0.235f
C732 ring_100mV_0.mdls_inv_3.OUT.n8 ss 0.235f
C733 ring_100mV_0.mdls_inv_3.OUT.n9 ss 0.306f
C734 ring_100mV_0.mdls_inv_3.OUT.t15 ss 0.255f
C735 ring_100mV_0.mdls_inv_3.OUT.t13 ss 0.255f
C736 ring_100mV_0.mdls_inv_3.OUT.t12 ss 0.255f
C737 ring_100mV_0.mdls_inv_3.OUT.t9 ss 0.255f
C738 ring_100mV_0.mdls_inv_3.OUT.t14 ss 0.374f
C739 ring_100mV_0.mdls_inv_3.OUT.n10 ss 0.393f
C740 ring_100mV_0.mdls_inv_3.OUT.t16 ss 0.255f
C741 ring_100mV_0.mdls_inv_3.OUT.n11 ss 0.238f
C742 ring_100mV_0.mdls_inv_3.OUT.n12 ss 0.238f
C743 ring_100mV_0.mdls_inv_3.OUT.t17 ss 0.255f
C744 ring_100mV_0.mdls_inv_3.OUT.n13 ss 0.238f
C745 ring_100mV_0.mdls_inv_3.OUT.n14 ss 0.238f
C746 ring_100mV_0.mdls_inv_3.OUT.t8 ss 0.255f
C747 ring_100mV_0.mdls_inv_3.OUT.n15 ss 0.238f
C748 ring_100mV_0.mdls_inv_3.OUT.n16 ss 0.224f
C749 ring_100mV_0.mdls_inv_3.OUT.n17 ss 0.151f
C750 ring_100mV_0.mdls_inv_3.OUT.n18 ss 0.529f
C751 ring_100mV_0.mdls_inv_3.OUT.t7 ss 0.118f
C752 ring_100mV_0.mdls_inv_3.OUT.t3 ss 0.00764f
C753 ring_100mV_0.mdls_inv_3.OUT.n19 ss 0.0878f
C754 ring_100mV_0.mdls_inv_3.OUT.n20 ss 0.225f
C755 ring_100mV_0.mdls_inv_3.OUT.n21 ss 0.319f
C756 ring_100mV_0.mdls_inv_3.OUT.t2 ss 0.465f
C757 ring_100mV_0.mdls_inv_3.OUT.t4 ss 0.465f
C758 ring_100mV_0.mdls_inv_3.OUT.t0 ss 0.496f
C759 ring_100mV_0.mdls_inv_3.OUT.n22 ss 0.138f
C760 ring_100mV_0.mdls_inv_3.OUT.n23 ss 0.133f
C761 ring_100mV_0.mdls_inv_3.OUT.t1 ss 0.042f
C762 ring_100mV_0.mdls_inv_3.OUT.n24 ss 0.35f
C763 iref_2nA_0.iref_2nA_mirrors_0.Ip1 ss 1.01f
C764 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t1 ss 0.0673f
C765 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t0 ss 0.0284f
C766 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t2 ss 0.0287f
C767 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t4 ss 0.591f
C768 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t6 ss 0.48f
C769 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n0 ss 1.69f
C770 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t5 ss 0.48f
C771 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n1 ss 0.904f
C772 iref_2nA_0.iref_2nA_igenerator_0.Ip1.t3 ss 0.48f
C773 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n2 ss 1.04f
C774 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n3 ss 0.889f
C775 iref_2nA_0.iref_2nA_igenerator_0.Ip1.n4 ss 0.765f
C776 ring_100mV_0.mdls_inv_6.IN.n0 ss 0.249f
C777 ring_100mV_0.mdls_inv_6.IN.n1 ss 0.261f
C778 ring_100mV_0.mdls_inv_6.IN.t11 ss 0.151f
C779 ring_100mV_0.mdls_inv_6.IN.t7 ss 0.151f
C780 ring_100mV_0.mdls_inv_6.IN.n2 ss 0.441f
C781 ring_100mV_0.mdls_inv_6.IN.t8 ss 0.194f
C782 ring_100mV_0.mdls_inv_6.IN.n3 ss 0.0758f
C783 ring_100mV_0.mdls_inv_6.IN.n4 ss 0.374f
C784 ring_100mV_0.mdls_inv_6.IN.n5 ss 0.484f
C785 ring_100mV_0.mdls_inv_6.IN.t6 ss 0.3f
C786 ring_100mV_0.mdls_inv_6.IN.t12 ss 0.298f
C787 ring_100mV_0.mdls_inv_6.IN.n6 ss 0.485f
C788 ring_100mV_0.mdls_inv_6.IN.t10 ss 0.299f
C789 ring_100mV_0.mdls_inv_6.IN.n7 ss 0.485f
C790 ring_100mV_0.mdls_inv_6.IN.t14 ss 0.298f
C791 ring_100mV_0.mdls_inv_6.IN.t13 ss 0.373f
C792 ring_100mV_0.mdls_inv_6.IN.n8 ss 0.293f
C793 ring_100mV_0.mdls_inv_6.IN.n9 ss 0.0975f
C794 ring_100mV_0.mdls_inv_6.IN.n10 ss 0.292f
C795 ring_100mV_0.mdls_inv_6.IN.t9 ss 0.373f
C796 ring_100mV_0.mdls_inv_6.IN.n11 ss 0.279f
C797 ring_100mV_0.mdls_inv_6.IN.t5 ss 0.402f
C798 ring_100mV_0.mdls_inv_6.IN.n12 ss 0.636f
C799 ring_100mV_0.mdls_inv_6.IN.n13 ss 0.594f
C800 ring_100mV_0.mdls_inv_6.IN.t15 ss 0.138f
C801 ring_100mV_0.mdls_inv_6.IN.t0 ss 0.00893f
C802 ring_100mV_0.mdls_inv_6.IN.n14 ss 0.103f
C803 ring_100mV_0.mdls_inv_6.IN.n15 ss 0.263f
C804 ring_100mV_0.mdls_inv_6.IN.n16 ss 0.373f
C805 ring_100mV_0.mdls_inv_6.IN.t2 ss 0.544f
C806 ring_100mV_0.mdls_inv_6.IN.t3 ss 0.58f
C807 ring_100mV_0.mdls_inv_6.IN.t1 ss 0.544f
C808 ring_100mV_0.mdls_inv_6.IN.n17 ss 0.162f
C809 ring_100mV_0.mdls_inv_6.IN.n18 ss 0.155f
C810 ring_100mV_0.mdls_inv_6.IN.t4 ss 0.0491f
C811 ring_100mV_0.mdls_inv_6.IN.n19 ss 0.409f
C812 ring_100mV_0.mdls_inv_8.OUT ss 0.0818f
C813 a_9754_13622.t2 ss 1.01f
C814 a_9754_13622.t4 ss 0.95f
C815 a_9754_13622.t1 ss 0.939f
C816 a_9754_13622.t3 ss 1.01f
C817 a_9754_13622.n0 ss 0.244f
C818 a_9754_13622.n1 ss 0.172f
C819 a_9754_13622.t6 ss 0.451f
C820 a_9754_13622.t0 ss 0.0858f
C821 a_9754_13622.n2 ss 0.91f
C822 a_9754_13622.n3 ss 0.154f
C823 a_9754_13622.n4 ss 0.234f
C824 a_9754_13622.t5 ss 0.946f
C825 dd_02.n0 ss 0.135f
C826 dd_02.n1 ss 0.118f
C827 dd_02.n2 ss 0.0083f
C828 dd_02.n3 ss 0.0656f
C829 dd_02.n4 ss 0.0656f
C830 dd_02.n5 ss 0.0656f
C831 ring_100mV_0.mdls_inv_1.DD ss 0.0185f
C832 dd_02.t18 ss 0.347f
C833 dd_02.t28 ss 0.337f
C834 dd_02.n6 ss 0.0985f
C835 dd_02.n7 ss 0.0424f
C836 dd_02.n8 ss 0.0487f
C837 dd_02.n9 ss 0.0656f
C838 dd_02.n10 ss 0.0487f
C839 dd_02.n11 ss 0.0656f
C840 dd_02.n12 ss 0.0487f
C841 dd_02.n13 ss 0.0656f
C842 dd_02.n14 ss 0.0487f
C843 dd_02.n15 ss 0.0656f
C844 dd_02.n16 ss 0.0487f
C845 dd_02.n17 ss 0.0653f
C846 dd_02.n18 ss 2.91f
C847 dd_02.t7 ss 0.347f
C848 dd_02.t4 ss 0.337f
C849 dd_02.n19 ss 0.0985f
C850 dd_02.n20 ss 0.0421f
C851 dd_02.n21 ss 0.0132f
C852 dd_02.n22 ss 0.0333f
C853 dd_02.n23 ss 2.16f
C854 dd_02.t5 ss 0.0683f
C855 dd_02.t35 ss 0.00529f
C856 dd_02.n24 ss 0.0902f
C857 dd_02.n25 ss 0.0311f
C858 dd_02.n26 ss 0.0661f
C859 dd_02.n27 ss 0.0665f
C860 dd_02.n28 ss 0.0665f
C861 dd_02.t31 ss 0.347f
C862 dd_02.t29 ss 0.337f
C863 dd_02.n29 ss 0.0985f
C864 dd_02.n30 ss 0.0424f
C865 dd_02.t32 ss 0.347f
C866 dd_02.t26 ss 0.337f
C867 dd_02.n31 ss 0.0985f
C868 dd_02.n32 ss 0.0424f
C869 dd_02.n33 ss 2.17f
C870 dd_02.n34 ss 0.0105f
C871 dd_02.n35 ss 0.0314f
C872 ring_100mV_0.mdls_inv_3.DD ss 0.0414f
C873 dd_02.n36 ss 0.00592f
C874 dd_02.n37 ss 0.00753f
C875 dd_02.t33 ss 0.00529f
C876 dd_02.n38 ss 0.0902f
C877 dd_02.n39 ss 0.0311f
C878 dd_02.n40 ss 0.0661f
C879 dd_02.t37 ss 0.347f
C880 dd_02.t39 ss 0.337f
C881 dd_02.n41 ss 0.0985f
C882 dd_02.n42 ss 0.0424f
C883 dd_02.n43 ss 0.0198f
C884 ring_100mV_0.mdls_inv_5.DD ss 0.0217f
C885 dd_02.n44 ss 0.136f
C886 dd_02.n45 ss 0.209f
C887 dd_02.n46 ss 0.131f
C888 ring_100mV_0.mdls_inv_4.DD ss 0.0185f
C889 dd_02.t34 ss 0.347f
C890 dd_02.t36 ss 0.337f
C891 dd_02.n47 ss 0.0985f
C892 dd_02.n48 ss 0.0424f
C893 dd_02.n49 ss 0.0189f
C894 dd_02.n50 ss 0.0665f
C895 dd_02.t14 ss 0.00529f
C896 dd_02.n51 ss 0.0902f
C897 dd_02.n52 ss 0.0311f
C898 dd_02.n53 ss 0.0665f
C899 dd_02.t10 ss 0.347f
C900 dd_02.t9 ss 0.337f
C901 dd_02.n54 ss 0.0985f
C902 dd_02.n55 ss 0.0424f
C903 dd_02.n56 ss 0.0198f
C904 ring_100mV_0.mdls_inv_7.DD ss 0.0217f
C905 dd_02.n57 ss 0.136f
C906 dd_02.n58 ss 0.209f
C907 dd_02.n59 ss 0.131f
C908 ring_100mV_0.mdls_inv_6.DD ss 0.0185f
C909 dd_02.t11 ss 0.347f
C910 dd_02.t12 ss 0.337f
C911 dd_02.n60 ss 0.0985f
C912 dd_02.n61 ss 0.0424f
C913 dd_02.n62 ss 0.0189f
C914 dd_02.n63 ss 0.0665f
C915 dd_02.t13 ss 0.00529f
C916 dd_02.n64 ss 0.0902f
C917 dd_02.n65 ss 0.0311f
C918 dd_02.n66 ss 0.0665f
C919 dd_02.t15 ss 0.00529f
C920 dd_02.n67 ss 0.0902f
C921 dd_02.n68 ss 0.0311f
C922 dd_02.n69 ss 0.0665f
C923 dd_02.t27 ss 0.347f
C924 dd_02.t19 ss 0.337f
C925 dd_02.n70 ss 0.0985f
C926 dd_02.n71 ss 0.0424f
C927 dd_02.n72 ss 0.0189f
C928 dd_02.n73 ss 0.0665f
C929 dd_02.n74 ss 0.0487f
C930 dd_02.n75 ss 0.0656f
C931 dd_02.n76 ss 0.0487f
C932 dd_02.n77 ss 0.0656f
C933 dd_02.n78 ss 0.0487f
C934 dd_02.n79 ss 0.0656f
C935 dd_02.n80 ss 0.0487f
C936 dd_02.n81 ss 0.0656f
C937 dd_02.n82 ss 0.0487f
C938 dd_02.n83 ss 0.0652f
C939 dd_02.n84 ss 2.88f
C940 dd_02.t40 ss 0.347f
C941 dd_02.t3 ss 0.337f
C942 dd_02.n85 ss 0.0985f
C943 dd_02.n86 ss 0.042f
C944 dd_02.n87 ss 0.0132f
C945 dd_02.n88 ss 0.0333f
C946 dd_02.n89 ss 2.16f
C947 dd_02.t2 ss 0.0911f
C948 dd_02.t43 ss 0.00529f
C949 dd_02.n90 ss 0.0902f
C950 dd_02.n91 ss 0.0311f
C951 dd_02.n92 ss 0.0665f
C952 dd_02.n93 ss 1.76f
C953 dd_02.n94 ss 0.0665f
C954 dd_02.n95 ss 0.0189f
C955 ring_100mV_0.mdls_inv_8.DD ss 0.0185f
C956 dd_02.n96 ss 0.136f
C957 dd_02.n97 ss 0.209f
C958 dd_02.n98 ss 0.131f
C959 ring_100mV_0.mdls_inv_9.DD ss 0.0217f
C960 dd_02.n99 ss 0.0198f
C961 dd_02.n100 ss 0.0665f
C962 dd_02.n101 ss 0.0656f
C963 dd_02.n102 ss 0.0656f
C964 dd_02.n103 ss 0.0656f
C965 dd_02.n104 ss 0.0656f
C966 dd_02.n105 ss 0.0228f
C967 dd_02.n106 ss 0.0328f
C968 dd_02.n108 ss 0.0228f
C969 dd_02.n109 ss 0.0109f
C970 dd_02.n110 ss 0.0281f
C971 dd_02.n111 ss 0.0106f
C972 dd_02.n112 ss 0.0593f
C973 ring_100mV_0.mdls_inv_2.DD ss 0.00537f
C974 dd_02.n113 ss 0.0194f
C975 dd_02.n115 ss 0.0405f
C976 dd_02.n116 ss 0.0258f
C977 dd_02.n117 ss 1.28f
C978 dd_02.n118 ss 2.17f
C979 dd_02.t30 ss 0.00529f
C980 dd_02.n119 ss 0.0902f
C981 dd_02.n120 ss 0.0311f
C982 dd_02.n121 ss 0.0665f
C983 dd_02.t8 ss 0.00529f
C984 dd_02.n122 ss 0.0902f
C985 dd_02.n123 ss 0.0311f
C986 dd_02.n124 ss 0.0665f
C987 dd_02.t38 ss 0.00529f
C988 dd_02.n125 ss 0.0902f
C989 dd_02.n126 ss 0.0311f
C990 dd_02.n127 ss 0.0665f
C991 dd_02.t6 ss 0.00529f
C992 dd_02.n128 ss 0.0902f
C993 dd_02.n129 ss 0.0311f
C994 dd_02.n130 ss 0.0665f
C995 dd_02.n131 ss 0.00642f
C996 dd_02.n132 ss 0.00753f
C997 dd_02.n133 ss 1.78f
C998 dd_02.n134 ss 0.0665f
C999 dd_02.n135 ss 0.0198f
C1000 dd_02.n136 ss 0.131f
C1001 dd_02.n137 ss 0.127f
C1002 dd_02.n138 ss 0.209f
C1003 dd_02.n139 ss 0.0656f
C1004 dd_02.n140 ss 0.0951f
C1005 dd_02.n141 ss 0.0228f
C1006 dd_02.n142 ss 0.134f
C1007 dd_02.n143 ss 0.107f
C1008 dd_02.n144 ss 0.0328f
C1009 dd_02.n146 ss 1.31f
C1010 dd_02.n147 ss 0.026f
C1011 dd_02.n148 ss 0.0435f
C1012 dd_02.n149 ss 0.0297f
C1013 dd_02.n150 ss 0.0239f
C1014 dd_02.n151 ss 0.238f
C1015 dd_02.t21 ss 0.00576f
C1016 dd_02.t23 ss 0.00576f
C1017 dd_02.n152 ss 0.114f
C1018 dd_02.t17 ss 0.0098f
C1019 dd_02.n153 ss 0.155f
C1020 dd_02.t25 ss 0.0097f
C1021 dd_02.n154 ss 0.148f
C1022 dd_02.n155 ss 0.061f
C1023 dd_02.n156 ss 0.127f
C1024 dd_02.n157 ss 0.0839f
C1025 dd_02.n158 ss 0.0838f
C1026 dd_02.n159 ss 0.0824f
C1027 dd_02.n160 ss 0.0842f
C1028 dd_02.n161 ss 0.081f
C1029 dd_02.n162 ss 0.547f
C1030 dd_02.t16 ss 0.668f
C1031 dd_02.t20 ss 0.547f
C1032 dd_02.n163 ss 0.364f
C1033 dd_02.t22 ss 0.545f
C1034 dd_02.t24 ss 0.668f
C1035 dd_02.t41 ss 0.518f
C1036 dd_02.n164 ss 0.0593f
C1037 dd_02.n165 ss 0.0593f
C1038 dd_02.n166 ss 0.114f
C1039 dd_02.t1 ss 0.0297f
C1040 dd_02.t42 ss 0.0295f
C1041 dd_02.n167 ss 0.0681f
C1042 dd_02.n168 ss 0.0593f
C1043 dd_02.n169 ss 0.364f
C1044 dd_02.t0 ss 0.518f
C1045 dd_02.n170 ss 0.543f
C1046 dd_02.n171 ss 0.059f
C1047 dd_02.n172 ss 0.0744f
C1048 dd_02.n173 ss 0.0291f
C1049 dd_02.n174 ss 0.0598f
C1050 dd_02.n175 ss 0.477f
C1051 dd_02.n176 ss 0.444f
C1052 dd_02.n177 ss 0.0847f
C1053 dd_02.n178 ss 0.0189f
C1054 dd_02.n179 ss 0.38f
C1055 ring_100mV_0.ring_100mV_buffer_0.DD ss 0.156f
C1056 dd_02.n180 ss 0.474f
C1057 ring_100mV_0.DD ss 1.94f
C1058 dd_01.t28 ss 0.0493f
C1059 dd_01.t21 ss 0.0423f
C1060 dd_01.n0 ss 0.189f
C1061 vref01_0.DD ss 0.0106f
C1062 dd_01.n1 ss 0.0301f
C1063 dd_01.n2 ss 0.357f
C1064 dd_01.n3 ss 0.0305f
C1065 dd_01.n4 ss 0.0305f
C1066 dd_01.t76 ss 0.509f
C1067 dd_01.n7 ss 0.0305f
C1068 dd_01.n8 ss 0.0226f
C1069 dd_01.n9 ss 0.358f
C1070 dd_01.n10 ss 0.0213f
C1071 dd_01.n11 ss 0.0556f
C1072 dd_01.n12 ss 0.878f
C1073 dd_01.n13 ss 0.0158f
C1074 dd_01.n14 ss 0.0178f
C1075 dd_01.t38 ss 0.00959f
C1076 dd_01.n16 ss 0.137f
C1077 dd_01.n17 ss 0.0185f
C1078 dd_01.n18 ss 0.0185f
C1079 dd_01.t37 ss 0.204f
C1080 dd_01.n20 ss 0.137f
C1081 dd_01.n21 ss 0.0185f
C1082 dd_01.n22 ss 0.0712f
C1083 dd_01.n23 ss 0.0989f
C1084 dd_01.n24 ss 0.272f
C1085 dd_01.n25 ss 0.222f
C1086 dd_01.t54 ss 0.17f
C1087 dd_01.n26 ss 0.0465f
C1088 dd_01.t67 ss 0.00782f
C1089 dd_01.n27 ss 0.0438f
C1090 dd_01.t64 ss 0.17f
C1091 dd_01.t57 ss 0.00782f
C1092 dd_01.n28 ss 0.0377f
C1093 dd_01.n29 ss 0.0263f
C1094 dd_01.n30 ss 0.0465f
C1095 dd_01.t55 ss 0.338f
C1096 dd_01.t74 ss 0.414f
C1097 dd_01.t26 ss 0.305f
C1098 dd_01.n31 ss 0.207f
C1099 dd_01.t35 ss 0.316f
C1100 dd_01.t29 ss 0.414f
C1101 dd_01.t65 ss 0.327f
C1102 dd_01.n32 ss 0.211f
C1103 dd_01.n33 ss 0.164f
C1104 dd_01.t66 ss 0.00165f
C1105 dd_01.n34 ss 0.0852f
C1106 dd_01.t30 ss 0.00165f
C1107 dd_01.n35 ss 0.0705f
C1108 dd_01.t36 ss 0.00165f
C1109 dd_01.n36 ss 0.0575f
C1110 dd_01.n37 ss 0.0277f
C1111 dd_01.t27 ss 0.00165f
C1112 dd_01.n38 ss 0.0559f
C1113 dd_01.t75 ss 0.00165f
C1114 dd_01.n39 ss 0.0705f
C1115 dd_01.t56 ss 0.00165f
C1116 dd_01.n40 ss 0.107f
C1117 dd_01.n41 ss 0.324f
C1118 dd_01.n42 ss 0.0842f
C1119 ldo_0.DD ss 0.938f
C1120 dd_01.n43 ss 3.44f
C1121 dd_01.n44 ss 6.29f
C1122 dd_01.t20 ss 0.00597f
C1123 dd_01.n45 ss 0.123f
C1124 dd_01.n46 ss 0.0302f
C1125 dd_01.t18 ss 0.39f
C1126 dd_01.n47 ss 0.194f
C1127 dd_01.n48 ss 0.0484f
C1128 dd_01.t19 ss 0.00464f
C1129 dd_01.n49 ss 0.0314f
C1130 dd_01.t59 ss 0.00379f
C1131 dd_01.t50 ss 0.00379f
C1132 dd_01.t6 ss 0.00464f
C1133 dd_01.n50 ss 0.115f
C1134 dd_01.t14 ss 0.00464f
C1135 dd_01.n51 ss 0.115f
C1136 dd_01.t11 ss 0.00464f
C1137 dd_01.n52 ss 0.105f
C1138 dd_01.t49 ss 9.28e-19
C1139 dd_01.n53 ss 0.0626f
C1140 dd_01.t48 ss 0.0724f
C1141 dd_01.n54 ss 0.061f
C1142 dd_01.n55 ss 0.0204f
C1143 dd_01.t63 ss 0.00379f
C1144 dd_01.t12 ss 0.00464f
C1145 dd_01.n56 ss 0.115f
C1146 dd_01.t16 ss 0.00464f
C1147 dd_01.n57 ss 0.115f
C1148 dd_01.t7 ss 0.00464f
C1149 dd_01.n58 ss 0.115f
C1150 dd_01.t10 ss 0.00464f
C1151 dd_01.n59 ss 0.105f
C1152 dd_01.t62 ss 9.28e-19
C1153 dd_01.n60 ss 0.0648f
C1154 dd_01.t61 ss 0.0724f
C1155 dd_01.n61 ss 0.0752f
C1156 dd_01.n62 ss 0.0269f
C1157 dd_01.t43 ss 0.00379f
C1158 dd_01.t44 ss 0.00379f
C1159 dd_01.t40 ss 9.28e-19
C1160 dd_01.n63 ss 0.0166f
C1161 dd_01.n64 ss 0.0415f
C1162 dd_01.t39 ss 0.0292f
C1163 dd_01.t41 ss 9.28e-19
C1164 dd_01.n65 ss 0.0166f
C1165 dd_01.t52 ss 9.28e-19
C1166 dd_01.n66 ss 0.0119f
C1167 dd_01.t53 ss 9.28e-19
C1168 dd_01.n67 ss 0.0119f
C1169 dd_01.n68 ss 0.0618f
C1170 dd_01.n69 ss 0.0415f
C1171 dd_01.t51 ss 0.0292f
C1172 dd_01.n70 ss 0.0642f
C1173 dd_01.n71 ss 0.0202f
C1174 dd_01.t22 ss 1.04f
C1175 dd_01.n72 ss 0.0457f
C1176 dd_01.n73 ss 0.866f
C1177 dd_01.t24 ss 1.04f
C1178 dd_01.t73 ss 9.28e-19
C1179 dd_01.n74 ss 0.0119f
C1180 dd_01.t72 ss 9.28e-19
C1181 dd_01.n75 ss 0.0119f
C1182 dd_01.n76 ss 0.148f
C1183 dd_01.n77 ss 0.022f
C1184 dd_01.n78 ss 0.0415f
C1185 dd_01.t71 ss 0.0292f
C1186 dd_01.n79 ss 0.0627f
C1187 dd_01.n80 ss 0.0234f
C1188 dd_01.t46 ss 9.28e-19
C1189 dd_01.n81 ss 0.0119f
C1190 dd_01.t47 ss 9.28e-19
C1191 dd_01.n82 ss 0.0119f
C1192 dd_01.n83 ss 0.0558f
C1193 dd_01.n84 ss 0.0415f
C1194 dd_01.t45 ss 0.0292f
C1195 dd_01.n85 ss 0.0627f
C1196 dd_01.n86 ss 0.0191f
C1197 dd_01.n87 ss 0.00795f
C1198 dd_01.n88 ss 0.0607f
C1199 dd_01.n89 ss 0.913f
C1200 dd_01.n90 ss 0.0607f
C1201 dd_01.n91 ss 0.0194f
C1202 dd_01.n92 ss 0.0861f
C1203 dd_01.t31 ss 0.0199f
C1204 dd_01.t25 ss 0.0199f
C1205 dd_01.t23 ss 0.0199f
C1206 dd_01.t32 ss 0.0199f
C1207 dd_01.n93 ss 0.152f
C1208 dd_01.n94 ss 0.117f
C1209 dd_01.n95 ss 1.3f
C1210 dd_01.n96 ss 0.0604f
C1211 dd_01.n97 ss 0.0652f
C1212 dd_01.n98 ss 0.115f
C1213 dd_01.n99 ss 0.149f
C1214 dd_01.n100 ss 0.102f
C1215 dd_01.n101 ss 0.0275f
C1216 dd_01.t42 ss 0.0724f
C1217 dd_01.n102 ss 0.0608f
C1218 dd_01.n103 ss 0.0265f
C1219 dd_01.n104 ss 0.0135f
C1220 dd_01.n105 ss 0.144f
C1221 dd_01.t5 ss 0.00464f
C1222 dd_01.n106 ss 0.115f
C1223 dd_01.t17 ss 0.00464f
C1224 dd_01.n107 ss 0.115f
C1225 dd_01.t15 ss 0.00464f
C1226 dd_01.n108 ss 0.0941f
C1227 dd_01.t8 ss 0.00464f
C1228 dd_01.n109 ss 0.115f
C1229 dd_01.t13 ss 0.00464f
C1230 dd_01.n110 ss 0.115f
C1231 dd_01.t4 ss 0.00464f
C1232 dd_01.n111 ss 0.115f
C1233 dd_01.t9 ss 0.00464f
C1234 dd_01.n112 ss 0.0953f
C1235 dd_01.n113 ss 0.0406f
C1236 dd_01.n114 ss 1.08f
C1237 dd_01.t3 ss 3.66f
C1238 dd_01.n115 ss 0.218f
C1239 dd_01.n116 ss 1.1f
C1240 dd_01.t0 ss 3.33f
C1241 dd_01.n117 ss 2.65f
C1242 dd_01.n118 ss 0.144f
C1243 dd_01.n119 ss 0.0079f
C1244 dd_01.n120 ss 0.0201f
C1245 dd_01.t58 ss 0.0724f
C1246 dd_01.n121 ss 0.0571f
C1247 dd_01.t60 ss 0.00109f
C1248 dd_01.n122 ss 0.0979f
C1249 dd_01.n123 ss 0.0159f
C1250 dd_01.n124 ss 0.0926f
C1251 dd_01.n125 ss 0.0149f
C1252 dd_01.n126 ss 0.0304f
C1253 dd_01.n127 ss 0.291f
C1254 dd_01.t1 ss 0.391f
C1255 dd_01.t68 ss 0.0858f
C1256 dd_01.t70 ss 9.28e-19
C1257 dd_01.n128 ss 0.16f
C1258 dd_01.n129 ss 0.0439f
C1259 dd_01.n130 ss 0.321f
C1260 dd_01.n131 ss 0.0251f
C1261 dd_01.t34 ss 0.0044f
C1262 dd_01.n132 ss 0.0754f
C1263 dd_01.n133 ss 0.266f
C1264 dd_01.n134 ss 0.0364f
C1265 dd_01.t69 ss 0.254f
C1266 dd_01.t33 ss 0.217f
C1267 dd_01.t2 ss 0.455f
C1268 dd_01.n135 ss 0.0298f
C1269 dd_01.n136 ss 0.0363f
C1270 dd_01.n137 ss 0.473f
C1271 dd_01.n138 ss 0.0362f
C1272 dd_01.n139 ss 0.0236f
C1273 dd_01.n140 ss 0.0144f
C1274 dd_01.n141 ss 0.05f
C1275 dd_01.n142 ss 0.229f
C1276 iref_2nA_0.iref_2nA_vref_0.DD ss 0.131f
C1277 dd_01.n143 ss 0.0898f
C1278 dd_01.n144 ss 0.175f
C1279 dd_01.n145 ss 0.026f
C1280 dd_01.n146 ss 0.383f
C1281 dd_01.n147 ss 0.0283f
C1282 dd_01.n148 ss 0.027f
C1283 dd_01.n149 ss 0.0266f
C1284 dd_01.n150 ss 0.0166f
C1285 dd_01.n152 ss 0.00693f
C1286 dd_01.n153 ss 0.0674f
C1287 dd_01.n154 ss 0.572f
C1288 iref_2nA_0.DD ss 5.47f
C1289 a_1555_7968.n0 ss 1.32f
C1290 a_1555_7968.t2 ss 0.0129f
C1291 a_1555_7968.t3 ss 0.412f
C1292 a_1555_7968.t1 ss 0.412f
C1293 a_1555_7968.t5 ss 0.0128f
C1294 a_1555_7968.t4 ss 0.0128f
C1295 a_1555_7968.t0 ss 0.0128f
C1296 iref_2nA_0.iref_2nA_mirrors_0.Ip2 ss 2.08f
C1297 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n0 ss 0.731f
C1298 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n1 ss 1.43f
C1299 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t7 ss 0.0478f
C1300 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t10 ss 0.0205f
C1301 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n2 ss 0.591f
C1302 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t9 ss 0.0205f
C1303 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t0 ss 0.0205f
C1304 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t3 ss 0.0478f
C1305 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n3 ss 0.591f
C1306 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t11 ss 0.0478f
C1307 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t1 ss 0.0205f
C1308 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n4 ss 0.591f
C1309 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t6 ss 0.0205f
C1310 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t2 ss 0.0205f
C1311 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t8 ss 0.0478f
C1312 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n5 ss 0.591f
C1313 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t19 ss 1.02f
C1314 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t22 ss 1.08f
C1315 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t13 ss 1.08f
C1316 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t17 ss 1.08f
C1317 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t24 ss 1.08f
C1318 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t12 ss 1.08f
C1319 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t14 ss 1.08f
C1320 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t20 ss 1.08f
C1321 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t25 ss 1.08f
C1322 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t16 ss 1.08f
C1323 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t21 ss 1.08f
C1324 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t23 ss 1.08f
C1325 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t15 ss 0.719f
C1326 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t18 ss 0.658f
C1327 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n6 ss 1.2f
C1328 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t4 ss 0.0296f
C1329 iref_2nA_0.iref_2nA_igenerator_0.Ip2.t5 ss 0.0429f
C1330 iref_2nA_0.iref_2nA_igenerator_0.Ip2.n7 ss 1.01f
.ends


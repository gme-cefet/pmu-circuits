magic
tech sky130A
magscale 1 2
timestamp 1695346156
<< nwell >>
rect -246 -1373 246 1373
<< pmos >>
rect -50 754 50 1154
rect -50 118 50 518
rect -50 -518 50 -118
rect -50 -1154 50 -754
<< pdiff >>
rect -108 1142 -50 1154
rect -108 766 -96 1142
rect -62 766 -50 1142
rect -108 754 -50 766
rect 50 1142 108 1154
rect 50 766 62 1142
rect 96 766 108 1142
rect 50 754 108 766
rect -108 506 -50 518
rect -108 130 -96 506
rect -62 130 -50 506
rect -108 118 -50 130
rect 50 506 108 518
rect 50 130 62 506
rect 96 130 108 506
rect 50 118 108 130
rect -108 -130 -50 -118
rect -108 -506 -96 -130
rect -62 -506 -50 -130
rect -108 -518 -50 -506
rect 50 -130 108 -118
rect 50 -506 62 -130
rect 96 -506 108 -130
rect 50 -518 108 -506
rect -108 -766 -50 -754
rect -108 -1142 -96 -766
rect -62 -1142 -50 -766
rect -108 -1154 -50 -1142
rect 50 -766 108 -754
rect 50 -1142 62 -766
rect 96 -1142 108 -766
rect 50 -1154 108 -1142
<< pdiffc >>
rect -96 766 -62 1142
rect 62 766 96 1142
rect -96 130 -62 506
rect 62 130 96 506
rect -96 -506 -62 -130
rect 62 -506 96 -130
rect -96 -1142 -62 -766
rect 62 -1142 96 -766
<< nsubdiff >>
rect -210 1303 -114 1337
rect 114 1303 210 1337
rect -210 1241 -176 1303
rect 176 1241 210 1303
rect -210 -1303 -176 -1241
rect 176 -1303 210 -1241
rect -210 -1337 -114 -1303
rect 114 -1337 210 -1303
<< nsubdiffcont >>
rect -114 1303 114 1337
rect -210 -1241 -176 1241
rect 176 -1241 210 1241
rect -114 -1337 114 -1303
<< poly >>
rect -50 1235 50 1251
rect -50 1201 -34 1235
rect 34 1201 50 1235
rect -50 1154 50 1201
rect -50 707 50 754
rect -50 673 -34 707
rect 34 673 50 707
rect -50 657 50 673
rect -50 599 50 615
rect -50 565 -34 599
rect 34 565 50 599
rect -50 518 50 565
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -565 50 -518
rect -50 -599 -34 -565
rect 34 -599 50 -565
rect -50 -615 50 -599
rect -50 -673 50 -657
rect -50 -707 -34 -673
rect 34 -707 50 -673
rect -50 -754 50 -707
rect -50 -1201 50 -1154
rect -50 -1235 -34 -1201
rect 34 -1235 50 -1201
rect -50 -1251 50 -1235
<< polycont >>
rect -34 1201 34 1235
rect -34 673 34 707
rect -34 565 34 599
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -599 34 -565
rect -34 -707 34 -673
rect -34 -1235 34 -1201
<< locali >>
rect -210 1303 -114 1337
rect 114 1303 210 1337
rect -210 1241 -176 1303
rect 176 1241 210 1303
rect -50 1201 -34 1235
rect 34 1201 50 1235
rect -96 1142 -62 1158
rect -96 750 -62 766
rect 62 1142 96 1158
rect 62 750 96 766
rect -50 673 -34 707
rect 34 673 50 707
rect -50 565 -34 599
rect 34 565 50 599
rect -96 506 -62 522
rect -96 114 -62 130
rect 62 506 96 522
rect 62 114 96 130
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -522 -62 -506
rect 62 -130 96 -114
rect 62 -522 96 -506
rect -50 -599 -34 -565
rect 34 -599 50 -565
rect -50 -707 -34 -673
rect 34 -707 50 -673
rect -96 -766 -62 -750
rect -96 -1158 -62 -1142
rect 62 -766 96 -750
rect 62 -1158 96 -1142
rect -50 -1235 -34 -1201
rect 34 -1235 50 -1201
rect -210 -1303 -176 -1241
rect 176 -1303 210 -1241
rect -210 -1337 -114 -1303
rect 114 -1337 210 -1303
<< viali >>
rect -34 1201 34 1235
rect -96 766 -62 1142
rect 62 766 96 1142
rect -34 673 34 707
rect -34 565 34 599
rect -96 130 -62 506
rect 62 130 96 506
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -506 -62 -130
rect 62 -506 96 -130
rect -34 -599 34 -565
rect -34 -707 34 -673
rect -96 -1142 -62 -766
rect 62 -1142 96 -766
rect -34 -1235 34 -1201
<< metal1 >>
rect -46 1235 46 1241
rect -46 1201 -34 1235
rect 34 1201 46 1235
rect -46 1195 46 1201
rect -102 1142 -56 1154
rect -102 766 -96 1142
rect -62 766 -56 1142
rect -102 754 -56 766
rect 56 1142 102 1154
rect 56 766 62 1142
rect 96 766 102 1142
rect 56 754 102 766
rect -46 707 46 713
rect -46 673 -34 707
rect 34 673 46 707
rect -46 667 46 673
rect -46 599 46 605
rect -46 565 -34 599
rect 34 565 46 599
rect -46 559 46 565
rect -102 506 -56 518
rect -102 130 -96 506
rect -62 130 -56 506
rect -102 118 -56 130
rect 56 506 102 518
rect 56 130 62 506
rect 96 130 102 506
rect 56 118 102 130
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -130 -56 -118
rect -102 -506 -96 -130
rect -62 -506 -56 -130
rect -102 -518 -56 -506
rect 56 -130 102 -118
rect 56 -506 62 -130
rect 96 -506 102 -130
rect 56 -518 102 -506
rect -46 -565 46 -559
rect -46 -599 -34 -565
rect 34 -599 46 -565
rect -46 -605 46 -599
rect -46 -673 46 -667
rect -46 -707 -34 -673
rect 34 -707 46 -673
rect -46 -713 46 -707
rect -102 -766 -56 -754
rect -102 -1142 -96 -766
rect -62 -1142 -56 -766
rect -102 -1154 -56 -1142
rect 56 -766 102 -754
rect 56 -1142 62 -766
rect 96 -1142 102 -766
rect 56 -1154 102 -1142
rect -46 -1201 46 -1195
rect -46 -1235 -34 -1201
rect 34 -1235 46 -1201
rect -46 -1241 46 -1235
<< properties >>
string FIXED_BBOX -193 -1320 193 1320
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.5 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1696350080
<< metal3 >>
rect -586 1512 586 1540
rect -586 -1512 502 1512
rect 566 -1512 586 1512
rect -586 -1540 586 -1512
<< via3 >>
rect 502 -1512 566 1512
<< mimcap >>
rect -546 1460 254 1500
rect -546 -1460 -506 1460
rect 214 -1460 254 1460
rect -546 -1500 254 -1460
<< mimcapcontact >>
rect -506 -1460 214 1460
<< metal4 >>
rect 486 1512 582 1528
rect -507 1460 215 1461
rect -507 -1460 -506 1460
rect 214 -1460 215 1460
rect -507 -1461 215 -1460
rect 486 -1512 502 1512
rect 566 -1512 582 1512
rect 486 -1528 582 -1512
<< properties >>
string FIXED_BBOX -586 -1540 294 1540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4 l 15 val 127.22 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1697054415
<< nwell >>
rect -1334 -3224 33 -1036
<< psubdiff >>
rect -1459 -962 -1435 -845
rect 1653 -962 1677 -845
<< nsubdiff >>
rect -1298 -1106 -1238 -1072
rect -63 -1106 -3 -1072
rect -1298 -1132 -1264 -1106
rect -1298 -3154 -1264 -3128
rect -37 -1132 -3 -1106
rect -37 -3154 -3 -3128
rect -1298 -3188 -1238 -3154
rect -63 -3188 -3 -3154
<< psubdiffcont >>
rect -1435 -962 1653 -845
<< nsubdiffcont >>
rect -1238 -1106 -63 -1072
rect -1298 -3128 -1264 -1132
rect -37 -3128 -3 -1132
rect -1238 -3188 -63 -3154
<< locali >>
rect -1451 -962 -1435 -845
rect 1653 -962 1669 -845
rect -1298 -1078 -1238 -1072
rect -1434 -1106 -1238 -1078
rect -63 -1106 -3 -1072
rect -1434 -1132 -1264 -1106
rect -1434 -2176 -1298 -1132
rect -922 -1192 -749 -1106
rect -283 -1199 -239 -1106
rect -37 -1132 -3 -1106
rect 528 -1128 680 -1120
rect 467 -1130 843 -1128
rect -1009 -2312 -970 -2148
rect -1009 -2353 -106 -2312
rect -1009 -3028 -970 -2353
rect -146 -3028 -106 -2353
rect -1298 -3154 -1264 -3128
rect 366 -1214 843 -1130
rect 366 -1225 530 -1214
rect 359 -1244 530 -1225
rect 677 -1227 843 -1214
rect 1030 -1222 1053 -962
rect 1124 -1222 1149 -962
rect 677 -1244 850 -1227
rect 359 -1256 469 -1244
rect 108 -2554 347 -2504
rect 108 -2731 150 -2554
rect 303 -2731 347 -2554
rect 359 -2678 444 -1256
rect 739 -1266 850 -1244
rect 1030 -1245 1149 -1222
rect 765 -2680 850 -1266
rect 1519 -1688 1599 -1280
rect 1519 -2324 1599 -1916
rect 108 -2763 347 -2731
rect 1519 -2960 1599 -2552
rect -37 -3154 -3 -3128
rect -1298 -3188 -1238 -3154
rect -63 -3188 -3 -3154
rect 1074 -3283 1229 -3263
rect 1074 -3367 1101 -3283
rect 1202 -3367 1229 -3283
rect 1074 -3385 1229 -3367
rect 1519 -3596 1599 -3188
<< viali >>
rect 1053 -962 1124 -938
rect 1053 -1222 1124 -962
rect 150 -2731 303 -2554
rect 1101 -3367 1202 -3283
<< metal1 >>
rect 1030 -938 1149 -914
rect -1200 -2258 -1158 -1280
rect -521 -1543 -486 -1236
rect -403 -1238 -316 -1182
rect -216 -1238 -129 -1182
rect 1030 -1222 1053 -938
rect 1124 -1208 1149 -938
rect 1124 -1222 1400 -1208
rect 1030 -1240 1400 -1222
rect 1030 -1245 1149 -1240
rect -523 -2258 -486 -1543
rect 1066 -1447 1135 -1245
rect 1066 -1504 1337 -1447
rect 1066 -1788 1135 -1504
rect 1377 -1788 1469 -1771
rect 1066 -1820 1469 -1788
rect -316 -2258 -216 -2086
rect -1200 -2295 -216 -2258
rect -316 -2422 -216 -2295
rect 1066 -2090 1135 -1820
rect 1377 -1833 1469 -1820
rect 1066 -2147 1334 -2090
rect 1066 -2423 1135 -2147
rect 1377 -2423 1469 -2407
rect 1066 -2455 1469 -2423
rect 108 -2554 347 -2504
rect 108 -2610 150 -2554
rect -138 -2731 150 -2610
rect 303 -2731 347 -2554
rect -138 -2763 347 -2731
rect 538 -2873 670 -2700
rect 1066 -2733 1135 -2455
rect 1377 -2469 1469 -2455
rect 1066 -2790 1334 -2733
rect 1066 -2873 1135 -2790
rect 538 -2930 1135 -2873
rect 1066 -3058 1135 -2930
rect 1377 -3058 1469 -3043
rect 1066 -3062 1469 -3058
rect -344 -3263 -210 -3080
rect 1066 -3090 1752 -3062
rect 1066 -3167 1135 -3090
rect 1321 -3103 1752 -3090
rect 1321 -3105 1469 -3103
rect 1321 -3192 1387 -3105
rect -344 -3283 1229 -3263
rect -344 -3367 1101 -3283
rect 1202 -3367 1229 -3283
rect -344 -3385 1229 -3367
rect 1709 -3636 1752 -3103
rect 1464 -3677 1752 -3636
use sky130_fd_pr__pfet_01v8_9XRXHT  sky130_fd_pr__pfet_01v8_9XRXHT_0
timestamp 1695345667
transform 0 1 -845 -1 0 -1670
box -532 -337 532 337
use sky130_fd_pr__pfet_01v8_lvt_AUUK23  sky130_fd_pr__pfet_01v8_lvt_AUUK23_0
timestamp 1695345667
transform 0 1 -266 -1 0 -1634
box -494 -150 494 150
use sky130_fd_pr__pfet_01v8_lvt_G4T6DY  sky130_fd_pr__pfet_01v8_lvt_G4T6DY_0
timestamp 1695346156
transform 0 1 604 -1 0 -1953
box -893 -307 893 307
use sky130_fd_pr__pfet_01v8_lvt_XRKP42  sky130_fd_pr__pfet_01v8_lvt_XRKP42_0
timestamp 1695345667
transform 0 1 -553 -1 0 -2751
box -371 -443 371 443
use sky130_fd_pr__pfet_01v8_PDY5CA  sky130_fd_pr__pfet_01v8_PDY5CA_0
timestamp 1695346156
transform -1 0 1423 0 -1 -2438
box -246 -1373 246 1373
<< labels >>
flabel locali 1540 -2134 1596 -2074 0 FreeSans 1600 0 0 0 VREF
flabel locali -1406 -1312 -1342 -1242 0 FreeSans 1600 0 0 0 DD
flabel metal1 1081 -1520 1118 -1449 0 FreeSans 1600 0 0 0 SS
<< end >>

* NGSPICE file created from iref_2nA_vref.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_lvt_G4T6DY w_n893_n307# a_n755_n88# a_697_n88# a_n697_n185#
X0 a_697_n88# a_n697_n185# a_n755_n88# w_n893_n307# sky130_fd_pr__pfet_01v8_lvt ad=0.255 pd=2.34 as=0.255 ps=2.34 w=0.88 l=6.97
.ends

.subckt sky130_fd_pr__pfet_01v8_9XRXHT w_n532_n337# a_n496_n237# a_438_n237# a_n438_n334#
X0 a_438_n237# a_n438_n334# a_n496_n237# w_n532_n337# sky130_fd_pr__pfet_01v8 ad=0.687 pd=5.32 as=0.687 ps=5.32 w=2.37 l=4.38
.ends

.subckt sky130_fd_pr__pfet_01v8_PDY5CA a_50_n1154# w_n246_n1373# a_n108_n518# a_n108_118#
+ a_n108_754# a_n50_21# a_n50_n615# a_50_118# a_50_754# a_n50_n1251# a_n108_n1154#
+ a_n50_657# a_50_n518#
X0 a_50_n1154# a_n50_n1251# a_n108_n1154# w_n246_n1373# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X1 a_50_118# a_n50_21# a_n108_118# w_n246_n1373# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2 a_50_n518# a_n50_n615# a_n108_n518# w_n246_n1373# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X3 a_50_754# a_n50_657# a_n108_754# w_n246_n1373# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_XRKP42 a_n335_n343# a_277_n343# a_n277_n440# w_n371_n443#
X0 a_277_n343# a_n277_n440# a_n335_n343# w_n371_n443# sky130_fd_pr__pfet_01v8_lvt ad=0.995 pd=7.44 as=0.995 ps=7.44 w=3.43 l=2.77
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_AUUK23 a_n458_n50# w_n494_n150# a_n400_n147# a_400_n50#
X0 a_400_n50# a_n400_n147# a_n458_n50# w_n494_n150# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
.ends


* Top level circuit iref_2nA_vref

Xsky130_fd_pr__pfet_01v8_lvt_G4T6DY_0 li_359_n2678# li_359_n2678# SS li_359_n2678#
+ sky130_fd_pr__pfet_01v8_lvt_G4T6DY
Xsky130_fd_pr__pfet_01v8_9XRXHT_0 DD DD li_359_n2678# m1_n1200_n2295# sky130_fd_pr__pfet_01v8_9XRXHT
Xsky130_fd_pr__pfet_01v8_PDY5CA_0 SS VREF VREF VREF VREF SS SS SS SS SS VREF SS SS
+ sky130_fd_pr__pfet_01v8_PDY5CA
Xsky130_fd_pr__pfet_01v8_lvt_XRKP42_0 m1_n1200_n2295# VREF li_359_n2678# DD sky130_fd_pr__pfet_01v8_lvt_XRKP42
Xsky130_fd_pr__pfet_01v8_lvt_AUUK23_0 DD DD DD m1_n1200_n2295# sky130_fd_pr__pfet_01v8_lvt_AUUK23
.end


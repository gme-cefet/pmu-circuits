magic
tech sky130A
magscale 1 2
timestamp 1698332137
<< locali >>
rect -1047 19784 18654 20384
rect -1047 19173 764 19784
rect 5507 19629 12606 19784
rect -1047 7299 -494 19173
rect 16247 17627 17282 19784
rect 16247 17621 16975 17627
rect 5453 16160 5849 16212
rect 5453 15676 6006 16160
rect 5453 15629 5849 15676
rect 11510 15672 11938 16174
rect 18219 8636 18315 8780
rect 14296 7365 14665 7386
rect -1047 7076 2091 7299
rect 5959 7076 12804 7245
rect 14296 7076 15868 7365
rect 18155 7076 18635 7446
rect -1047 6476 18788 7076
rect -1047 6466 -494 6476
<< metal1 >>
rect 11103 17945 12417 17992
rect 11103 17720 11162 17945
rect 12344 17720 12417 17945
rect 11103 17676 12417 17720
rect 13052 16088 13638 20761
rect 15556 18292 18647 18571
rect 15556 17556 15835 18292
rect 15556 17552 15918 17556
rect 15556 17461 15931 17552
rect 15737 17423 15931 17461
rect 15798 17362 15931 17423
rect 12650 15851 13638 16088
rect 18368 15242 18647 18292
rect 16133 14963 18647 15242
rect 16133 14550 16412 14963
rect 13596 14124 18558 14550
rect 13597 13888 18558 14124
rect 13597 13886 18539 13888
rect 13599 13882 16256 13886
rect 4766 9676 5354 9772
rect 4766 7246 4854 9676
rect 5270 7246 5354 9676
rect 4766 7166 5354 7246
rect 4766 6140 5352 7166
rect 13599 6140 14090 13882
rect 17989 13735 18511 13886
rect 18067 10565 18686 10994
rect 18401 10009 18782 10214
rect 16311 7296 16465 7327
rect 16311 7117 18938 7296
rect -726 5482 18815 6140
<< via1 >>
rect 11162 17720 12344 17945
rect 4854 7246 5270 9676
<< metal2 >>
rect 12233 17992 12413 20748
rect 11103 17945 12417 17992
rect 11103 17720 11162 17945
rect 12344 17720 12417 17945
rect 11103 17676 12417 17720
rect 16482 15937 16626 16160
rect 16482 15844 18576 15937
rect 16483 15706 18576 15844
rect 4766 9676 5354 9760
rect 4766 7781 4854 9676
rect 4456 7246 4854 7781
rect 5270 7246 5354 9676
rect 4456 7243 5354 7246
rect 4766 7166 5354 7243
<< metal3 >>
rect -1074 8423 461 9174
rect 18391 8894 18870 9125
use iref_2nA  iref_2nA_0
timestamp 1698328096
transform 0 1 4468 -1 0 16274
box -3409 -5056 9048 205
use ldo  ldo_0
timestamp 1698328593
transform 1 0 5724 0 1 17576
box 8574 -10258 12913 -3712
use ring_100mV  ring_100mV_0
timestamp 1697065484
transform 1 0 4604 0 1 12805
box 848 -5593 8961 6935
use vref01  vref01_0
timestamp 1698329069
transform 1 0 16504 0 1 15556
box -2152 -116 1826 2666
<< labels >>
flabel metal2 12262 20580 12382 20694 0 FreeSans 3200 90 0 0 ring_out
port 0 nsew
flabel metal1 13290 20582 13410 20696 0 FreeSans 3200 90 0 0 dd_02
port 1 nsew
flabel metal2 17886 15766 18006 15880 0 FreeSans 3200 0 0 0 vref
port 2 nsew
flabel metal1 18374 10724 18494 10838 0 FreeSans 3200 0 0 0 ldo_out
port 3 nsew
flabel metal1 18674 10062 18748 10150 0 FreeSans 3200 0 0 0 ldo_vs
port 4 nsew
flabel metal3 18678 8958 18752 9046 0 FreeSans 3200 0 0 0 ldo_vb
port 5 nsew
flabel metal1 18716 7170 18790 7258 0 FreeSans 3200 0 0 0 ldo_iref
port 6 nsew
flabel metal1 18374 5776 18448 5864 0 FreeSans 3200 0 0 0 dd_01
port 7 nsew
flabel locali -718 6724 -526 6906 0 FreeSans 3200 0 0 0 ss
port 8 nsew
flabel metal3 -840 8674 -648 8856 0 FreeSans 3200 0 0 0 iref
port 9 nsew
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1697059911
<< locali >>
rect -1047 19784 18654 20384
rect -1047 7299 -494 19784
rect 5507 19629 12606 19784
rect 16247 17627 17282 19784
rect 16247 17621 16975 17627
rect 11510 15672 11938 16174
rect -1047 7076 2091 7299
rect 5959 7076 12804 7245
rect 14590 7076 15868 7365
rect -1047 6476 18788 7076
rect -1047 6466 -494 6476
<< metal1 >>
rect 11103 17945 12417 17992
rect 11103 17720 11162 17945
rect 12344 17720 12417 17945
rect 11103 17676 12417 17720
rect 13052 16088 13638 20761
rect 12650 15851 13638 16088
rect 14120 16972 15762 17227
rect 14120 14470 14593 16972
rect 13599 14255 14593 14470
rect 13597 13886 18539 14255
rect 4766 9676 5354 9772
rect 4766 7246 4854 9676
rect 5270 7246 5354 9676
rect 4766 7166 5354 7246
rect 4766 6140 5352 7166
rect 13599 6140 14090 13886
rect 17989 13735 18511 13886
rect 18067 10565 18686 10994
rect 18401 10009 18782 10214
rect 16311 7296 16465 7327
rect 16311 7117 18938 7296
rect -726 5482 18815 6140
<< via1 >>
rect 11162 17720 12344 17945
rect 4854 7246 5270 9676
<< metal2 >>
rect 12233 17992 12413 20748
rect 11103 17945 12417 17992
rect 11103 17720 11162 17945
rect 12344 17720 12417 17945
rect 11103 17676 12417 17720
rect 16482 15937 16626 16160
rect 16482 15844 18576 15937
rect 16483 15706 18576 15844
rect 4766 9676 5354 9760
rect 4766 7781 4854 9676
rect 4456 7246 4854 7781
rect 5270 7246 5354 9676
rect 4456 7243 5354 7246
rect 4766 7166 5354 7243
<< metal3 >>
rect -1074 8423 461 9174
rect 18391 8894 18870 9125
use iref_2nA  iref_2nA_0
timestamp 1697059543
transform 0 1 4468 -1 0 16274
box -3409 -5056 9048 205
use ldo  ldo_0
timestamp 1696513288
transform 1 0 5724 0 1 17576
box 8574 -10258 12913 -3712
use ring_100mV  ring_100mV_0
timestamp 1697040310
transform 1 0 4604 0 1 12805
box 848 -5593 8961 6935
use vref01  vref01_0
timestamp 1697049024
transform 1 0 16504 0 1 15556
box -1468 426 1392 2102
<< labels >>
flabel metal2 12268 20576 12374 20692 0 FreeSans 3200 90 0 0 ring_out
port 0 nsew
flabel metal1 13284 20576 13390 20692 0 FreeSans 3200 90 0 0 dd_02
port 1 nsew
flabel metal2 18374 15766 18480 15882 0 FreeSans 3200 0 0 0 vref
port 2 nsew
flabel metal1 18410 10834 18516 10950 0 FreeSans 3200 0 0 0 ldo_out
port 3 nsew
flabel metal1 18450 10064 18556 10180 0 FreeSans 3200 0 0 0 ldo_vs
port 4 nsew
flabel metal3 18678 8944 18784 9060 0 FreeSans 3200 0 0 0 ldo_vb
port 5 nsew
flabel metal1 18736 7148 18842 7264 0 FreeSans 3200 0 0 0 ldo_iref
port 6 nsew
flabel metal1 18338 5744 18444 5860 0 FreeSans 3200 0 0 0 dd_01
port 7 nsew
flabel metal3 -892 8714 -786 8830 0 FreeSans 3200 0 0 0 iref
port 8 nsew
flabel locali -854 6722 -748 6838 0 FreeSans 3200 0 0 0 ss
port 9 nsew
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1695828444
<< psubdiff >>
rect 3771 -1602 3926 -1529
rect 6324 -1602 6523 -1529
rect 3771 -1605 3859 -1602
rect 3771 -2368 3859 -2280
rect 3769 -2470 3859 -2368
rect 6435 -1621 6523 -1602
rect 3769 -2546 3793 -2470
rect 4423 -2546 4516 -2470
rect 6435 -2472 6523 -2296
rect 5815 -2566 5927 -2472
rect 6533 -2566 6557 -2472
<< psubdiffcont >>
rect 3926 -1602 6324 -1529
rect 3771 -2280 3859 -1605
rect 6435 -2296 6523 -1621
rect 3793 -2546 4423 -2470
rect 5927 -2566 6533 -2472
<< locali >>
rect 3771 -1605 3859 -1589
rect 3910 -1602 3926 -1529
rect 6324 -1602 6340 -1529
rect 3770 -2280 3771 -2266
rect 6435 -1621 6523 -1605
rect 3859 -1758 4267 -1686
rect 6020 -1758 6435 -1686
rect 4232 -2266 4267 -1758
rect 3859 -2280 4267 -2266
rect 3770 -2338 4267 -2280
rect 4232 -2376 4267 -2338
rect 3777 -2546 3793 -2470
rect 4423 -2546 4439 -2470
rect 4648 -2492 4683 -1758
rect 5064 -2371 5099 -1758
rect 5063 -2383 5099 -2371
rect 5480 -2383 5515 -1758
rect 5063 -2392 5515 -2383
rect 5063 -2421 5236 -2392
rect 5206 -2429 5236 -2421
rect 5356 -2421 5515 -2392
rect 5356 -2429 5379 -2421
rect 5206 -2436 5379 -2429
rect 5896 -2472 5931 -1758
rect 6312 -2266 6347 -1758
rect 6020 -2296 6435 -2266
rect 6020 -2338 6523 -2296
rect 6312 -2376 6347 -2338
rect 5811 -2521 5927 -2472
rect 5911 -2566 5927 -2521
rect 6533 -2566 6549 -2472
rect 5684 -2800 5807 -2699
<< viali >>
rect 5236 -2429 5356 -2392
<< metal1 >>
rect 4311 -1379 4464 -1355
rect 4311 -1435 4349 -1379
rect 4426 -1435 4464 -1379
rect 4311 -1452 4464 -1435
rect 4311 -2028 4361 -1452
rect 4727 -1461 5193 -1372
rect 5456 -1379 5609 -1355
rect 5456 -1435 5494 -1379
rect 5571 -1435 5609 -1379
rect 5456 -1452 5609 -1435
rect 4727 -2028 4777 -1461
rect 5143 -2028 5193 -1461
rect 5559 -2028 5609 -1452
rect 3990 -2340 4186 -2294
rect 4406 -2340 5846 -2294
rect 6066 -2340 6262 -2294
rect 5710 -2381 5809 -2340
rect 6574 -2381 6630 -1427
rect 5206 -2392 5379 -2385
rect 5206 -2402 5236 -2392
rect 4415 -2429 5236 -2402
rect 5356 -2429 5379 -2392
rect 4415 -2436 5379 -2429
rect 5710 -2431 6630 -2381
rect 4415 -2438 5333 -2436
rect 4415 -2749 4455 -2438
rect 5588 -2558 5857 -2535
rect 5588 -2568 6075 -2558
rect 4415 -2791 4630 -2749
rect 5825 -2924 6075 -2568
rect 5590 -2927 6075 -2924
rect 5590 -2957 5857 -2927
<< via1 >>
rect 4349 -1435 4426 -1379
rect 5494 -1435 5571 -1379
<< metal2 >>
rect 4311 -1379 4464 -1355
rect 4311 -1435 4349 -1379
rect 4426 -1386 4464 -1379
rect 5456 -1379 5609 -1355
rect 5456 -1386 5494 -1379
rect 4426 -1433 5494 -1386
rect 4426 -1435 4464 -1433
rect 4311 -1452 4464 -1435
rect 5456 -1435 5494 -1433
rect 5571 -1435 5609 -1379
rect 5456 -1452 5609 -1435
use sky130_fd_pr__nfet_01v8_lvt_4HNDKD  sky130_fd_pr__nfet_01v8_lvt_4HNDKD_0
timestamp 1695826972
transform 1 0 5161 0 1 -2746
box -696 -310 696 310
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_0
timestamp 1695788690
transform 1 0 4502 0 1 -2012
box -158 -338 158 338
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_1
timestamp 1695788690
transform 1 0 4086 0 1 -2012
box -158 -338 158 338
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_3
timestamp 1695788690
transform 1 0 5334 0 1 -2012
box -158 -338 158 338
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_4
timestamp 1695788690
transform 1 0 4918 0 1 -2012
box -158 -338 158 338
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_6
timestamp 1695788690
transform 1 0 5750 0 1 -2012
box -158 -338 158 338
use sky130_fd_pr__nfet_01v8_lvt_C9VRMX  sky130_fd_pr__nfet_01v8_lvt_C9VRMX_7
timestamp 1695788690
transform 1 0 6166 0 1 -2012
box -158 -338 158 338
<< labels >>
rlabel metal1 6580 -1498 6622 -1440 3 Vg
rlabel metal1 5146 -1690 5188 -1632 3 Ip1
rlabel metal1 5560 -1690 5602 -1632 3 Ip2
rlabel locali 5728 -2776 5770 -2718 3 SS
rlabel metal1 5932 -2796 5974 -2738 3 VCTAT
<< end >>

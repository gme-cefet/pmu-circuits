magic
tech sky130A
magscale 1 2
timestamp 1696347688
<< metal3 >>
rect -966 792 966 820
rect -966 -792 882 792
rect 946 -792 966 792
rect -966 -820 966 -792
<< via3 >>
rect 882 -792 946 792
<< mimcap >>
rect -926 740 634 780
rect -926 -740 -886 740
rect 594 -740 634 740
rect -926 -780 634 -740
<< mimcapcontact >>
rect -886 -740 594 740
<< metal4 >>
rect 866 792 962 808
rect -887 740 595 741
rect -887 -740 -886 740
rect 594 -740 595 740
rect -887 -741 595 -740
rect 866 -792 882 792
rect 946 -792 962 792
rect 866 -808 962 -792
<< properties >>
string FIXED_BBOX -966 -820 674 820
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 7.8 l 7.8 val 127.607 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1695405779
<< nwell >>
rect -294 -350 294 350
<< pmoslvt >>
rect -200 -250 200 250
<< pdiff >>
rect -258 238 -200 250
rect -258 -238 -246 238
rect -212 -238 -200 238
rect -258 -250 -200 -238
rect 200 238 258 250
rect 200 -238 212 238
rect 246 -238 258 238
rect 200 -250 258 -238
<< pdiffc >>
rect -246 -238 -212 238
rect 212 -238 246 238
<< poly >>
rect -200 331 200 347
rect -200 297 -184 331
rect 184 297 200 331
rect -200 250 200 297
rect -200 -297 200 -250
rect -200 -331 -184 -297
rect 184 -331 200 -297
rect -200 -347 200 -331
<< polycont >>
rect -184 297 184 331
rect -184 -331 184 -297
<< locali >>
rect -200 297 -184 331
rect 184 297 200 331
rect -246 238 -212 254
rect -246 -254 -212 -238
rect 212 238 246 254
rect 212 -254 246 -238
rect -200 -331 -184 -297
rect 184 -331 200 -297
<< viali >>
rect -184 297 184 331
rect -246 -238 -212 238
rect 212 -238 246 238
rect -184 -331 184 -297
<< metal1 >>
rect -196 331 196 337
rect -196 297 -184 331
rect 184 297 196 331
rect -196 291 196 297
rect -252 238 -206 250
rect -252 -238 -246 238
rect -212 -238 -206 238
rect -252 -250 -206 -238
rect 206 238 252 250
rect 206 -238 212 238
rect 246 -238 252 238
rect 206 -250 252 -238
rect -196 -297 196 -291
rect -196 -331 -184 -297
rect 184 -331 196 -297
rect -196 -337 196 -331
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2.5 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1697230679
use iref_2nA  iref_2nA_0
timestamp 1697064583
transform 0 1 4468 -1 0 16274
box -3409 -5056 9048 205
use ldo  ldo_0
timestamp 1697064844
transform 1 0 5724 0 1 17576
box 8574 -10258 12913 -3712
use ring_100mV  ring_100mV_0
timestamp 1697065484
transform 1 0 4604 0 1 12805
box 848 -5593 8961 6935
use vref01  vref01_0
timestamp 1697065228
transform 1 0 16504 0 1 15556
box -1468 426 1392 2102
<< end >>

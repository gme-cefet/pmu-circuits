magic
tech sky130A
timestamp 1695675331
<< error_p >>
rect -18 311 18 314
rect -18 294 -12 311
rect -18 291 18 294
rect -18 -294 18 -291
rect -18 -311 -12 -294
rect -18 -314 18 -311
<< nmoslvt >>
rect -20 -275 20 275
<< ndiff >>
rect -49 269 -20 275
rect -49 -269 -43 269
rect -26 -269 -20 269
rect -49 -275 -20 -269
rect 20 269 49 275
rect 20 -269 26 269
rect 43 -269 49 269
rect 20 -275 49 -269
<< ndiffc >>
rect -43 -269 -26 269
rect 26 -269 43 269
<< poly >>
rect -20 311 20 319
rect -20 294 -12 311
rect 12 294 20 311
rect -20 275 20 294
rect -20 -294 20 -275
rect -20 -311 -12 -294
rect 12 -311 20 -294
rect -20 -319 20 -311
<< polycont >>
rect -12 294 12 311
rect -12 -311 12 -294
<< locali >>
rect -20 294 -12 311
rect 12 294 20 311
rect -43 269 -26 277
rect -43 -277 -26 -269
rect 26 269 43 277
rect 26 -277 43 -269
rect -20 -311 -12 -294
rect 12 -311 20 -294
<< viali >>
rect -12 294 12 311
rect -43 -269 -26 269
rect 26 -269 43 269
rect -12 -311 12 -294
<< metal1 >>
rect -18 311 18 314
rect -18 294 -12 311
rect 12 294 18 311
rect -18 291 18 294
rect -46 269 -23 275
rect -46 -269 -43 269
rect -26 -269 -23 269
rect -46 -275 -23 -269
rect 23 269 46 275
rect 23 -269 26 269
rect 43 -269 46 269
rect 23 -275 46 -269
rect -18 -294 18 -291
rect -18 -311 -12 -294
rect 12 -311 18 -294
rect -18 -314 18 -311
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.5 l 0.4 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_lvt_5VYM7K a_n66_n598# a_n124_n510# a_66_n510# VSUBS
X0 a_66_n510# a_n66_n598# a_n124_n510# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
.ends

.subckt sky130_fd_pr__pfet_01v8_TRB9BZ a_n389_n186# w_n483_n189# a_n447_n89# a_389_n89#
X0 a_389_n89# a_n389_n186# a_n447_n89# w_n483_n189# sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_8D4JM4 a_n127_n704# w_n221_n707# a_n185_n607#
+ a_127_n607#
X0 a_127_n607# a_n127_n704# a_n185_n607# w_n221_n707# sky130_fd_pr__pfet_01v8_lvt ad=1.76 pd=12.7 as=1.76 ps=12.7 w=6.07 l=1.27
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_4FSB7X c1_n546_n1500# m3_n586_n1540#
X0 c1_n546_n1500# m3_n586_n1540# sky130_fd_pr__cap_mim_m3_1 l=15 w=4
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_EFQJD4 a_n95_n517# a_37_n517# a_n37_n614# w_n233_n736#
X0 a_37_n517# a_n37_n614# a_n95_n517# w_n233_n736# sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.9 as=1.5 ps=10.9 w=5.17 l=0.37
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_W6ELF5 a_n143_n1235# a_n201_109# a_143_n1147#
+ a_143_109# a_n143_21# a_n201_n1147# a_n303_n1321#
X0 a_143_n1147# a_n143_n1235# a_n201_n1147# a_n303_n1321# sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=5.19 l=1.43
X1 a_143_109# a_n143_21# a_n201_109# a_n303_n1321# sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=5.19 l=1.43
.ends

.subckt ldo Iref SS VB VS OUT DD
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_0 Iref Iref SS SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_1 SS SS SS SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_2 Iref SS m1_9175_n5154# SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_3 Iref SS m1_9116_n8088# SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_5 Iref SS Iref SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_4 Iref SS m1_9116_n8088# SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_6 Iref m1_9116_n8088# SS SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__pfet_01v8_TRB9BZ_0 DD DD DD DD sky130_fd_pr__pfet_01v8_TRB9BZ
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_7 Iref m1_9116_n8088# SS SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_8 SS SS SS SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__pfet_01v8_TRB9BZ_2 m1_9175_n5154# DD DD m1_8616_n5605# sky130_fd_pr__pfet_01v8_TRB9BZ
Xsky130_fd_pr__pfet_01v8_TRB9BZ_1 DD DD DD DD sky130_fd_pr__pfet_01v8_TRB9BZ
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_9 Iref m1_9175_n5154# SS SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__pfet_01v8_TRB9BZ_3 m1_9175_n5154# DD DD m1_9175_n5154# sky130_fd_pr__pfet_01v8_TRB9BZ
Xsky130_fd_pr__pfet_01v8_TRB9BZ_4 m1_9175_n5154# DD DD m1_9175_n5154# sky130_fd_pr__pfet_01v8_TRB9BZ
Xsky130_fd_pr__pfet_01v8_TRB9BZ_5 m1_9175_n5154# DD DD m1_8616_n5605# sky130_fd_pr__pfet_01v8_TRB9BZ
Xsky130_fd_pr__pfet_01v8_lvt_8D4JM4_0 VS OUT OUT m1_9116_n8088# sky130_fd_pr__pfet_01v8_lvt_8D4JM4
Xsky130_fd_pr__pfet_01v8_lvt_8D4JM4_1 VS OUT OUT m1_9116_n8088# sky130_fd_pr__pfet_01v8_lvt_8D4JM4
Xsky130_fd_pr__cap_mim_m3_1_4FSB7X_0 m1_8616_n5605# OUT sky130_fd_pr__cap_mim_m3_1_4FSB7X
Xsky130_fd_pr__pfet_01v8_lvt_EFQJD4_0 DD OUT m1_8616_n5605# DD sky130_fd_pr__pfet_01v8_lvt_EFQJD4
Xsky130_fd_pr__nfet_01v8_lvt_W6ELF5_0 VB m1_8616_n5605# m1_9116_n8088# m1_9116_n8088#
+ VB m1_8616_n5605# SS sky130_fd_pr__nfet_01v8_lvt_W6ELF5
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_62AYNZ a_n158_n550# a_n100_n638# a_100_n550# VSUBS
X0 a_100_n550# a_n100_n638# a_n158_n550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_P9XYHJ a_80_n550# a_n138_n550# a_n80_n638# VSUBS
X0 a_80_n550# a_n80_n638# a_n138_n550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.8
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_G2G9KE a_n138_n100# a_n80_n197# a_80_n100# w_n174_n200#
X0 a_80_n100# a_n80_n197# a_n138_n100# w_n174_n200# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.8
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_NCVK88 a_n258_n100# a_n200_n197# a_200_n100# w_n294_n200#
X0 a_200_n100# a_n200_n197# a_n258_n100# w_n294_n200# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_P34KHJ a_40_n550# a_n98_n550# a_n40_n638# VSUBS
X0 a_40_n550# a_n40_n638# a_n98_n550# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.4
.ends

.subckt mdls_inv a_2701_260# OUT IN DD SS
Xsky130_fd_pr__nfet_01v8_lvt_62AYNZ_1 li_n14_266# IN SS SS sky130_fd_pr__nfet_01v8_lvt_62AYNZ
Xsky130_fd_pr__nfet_01v8_lvt_62AYNZ_0 li_n14_266# IN SS SS sky130_fd_pr__nfet_01v8_lvt_62AYNZ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_4 OUT li_n14_266# IN SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_5 OUT li_n14_266# IN SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_6 OUT li_n14_266# IN SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_7 OUT li_n14_266# IN SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__pfet_01v8_lvt_G2G9KE_0 m1_2309_1084# IN OUT DD sky130_fd_pr__pfet_01v8_lvt_G2G9KE
Xsky130_fd_pr__pfet_01v8_lvt_G2G9KE_1 li_n14_266# OUT SS DD sky130_fd_pr__pfet_01v8_lvt_G2G9KE
Xsky130_fd_pr__pfet_01v8_lvt_NCVK88_0 m1_2309_1084# IN DD DD sky130_fd_pr__pfet_01v8_lvt_NCVK88
Xsky130_fd_pr__nfet_01v8_lvt_P34KHJ_0 m1_2309_1084# DD OUT SS sky130_fd_pr__nfet_01v8_lvt_P34KHJ
Xsky130_fd_pr__nfet_01v8_lvt_P34KHJ_1 m1_2309_1084# DD OUT SS sky130_fd_pr__nfet_01v8_lvt_P34KHJ
.ends

.subckt ring_100mV_buffer OUT IN DD SS
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_28 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_29 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_0 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_17 SS li_8388_n2876# IN SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_18 SS li_8388_n2876# IN SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_1 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_19 SS li_8388_n2876# IN SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_2 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_3 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_4 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_5 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_6 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_7 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_8 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__pfet_01v8_lvt_G2G9KE_0 li_8388_n2876# IN DD DD sky130_fd_pr__pfet_01v8_lvt_G2G9KE
Xsky130_fd_pr__pfet_01v8_lvt_G2G9KE_1 DD IN li_8388_n2876# DD sky130_fd_pr__pfet_01v8_lvt_G2G9KE
Xsky130_fd_pr__pfet_01v8_lvt_G2G9KE_2 DD li_8388_n2876# OUT DD sky130_fd_pr__pfet_01v8_lvt_G2G9KE
Xsky130_fd_pr__pfet_01v8_lvt_G2G9KE_3 OUT li_8388_n2876# DD DD sky130_fd_pr__pfet_01v8_lvt_G2G9KE
Xsky130_fd_pr__pfet_01v8_lvt_G2G9KE_4 OUT li_8388_n2876# DD DD sky130_fd_pr__pfet_01v8_lvt_G2G9KE
Xsky130_fd_pr__pfet_01v8_lvt_G2G9KE_5 DD li_8388_n2876# OUT DD sky130_fd_pr__pfet_01v8_lvt_G2G9KE
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_30 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_31 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_20 SS li_8388_n2876# IN SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_21 SS li_8388_n2876# IN SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_22 SS li_8388_n2876# IN SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_23 SS li_8388_n2876# IN SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_25 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_26 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_27 OUT SS li_8388_n2876# SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
Xsky130_fd_pr__nfet_01v8_lvt_P9XYHJ_16 SS li_8388_n2876# IN SS sky130_fd_pr__nfet_01v8_lvt_P9XYHJ
.ends

.subckt ring_100mV SS DD ring_100mV_buffer_0/OUT
Xmdls_inv_0 SS mdls_inv_1/IN mdls_inv_0/IN DD SS mdls_inv
Xmdls_inv_1 SS mdls_inv_8/IN mdls_inv_1/IN DD SS mdls_inv
Xmdls_inv_2 SS mdls_inv_5/IN mdls_inv_3/IN DD SS mdls_inv
Xmdls_inv_3 SS mdls_inv_3/OUT mdls_inv_3/IN DD SS mdls_inv
Xmdls_inv_4 SS mdls_inv_3/IN mdls_inv_4/IN DD SS mdls_inv
Xmdls_inv_5 SS mdls_inv_7/IN mdls_inv_5/IN DD SS mdls_inv
Xmdls_inv_6 SS mdls_inv_4/IN mdls_inv_6/IN DD SS mdls_inv
Xmdls_inv_7 SS mdls_inv_9/IN mdls_inv_7/IN DD SS mdls_inv
Xmdls_inv_9 SS mdls_inv_0/IN mdls_inv_9/IN DD SS mdls_inv
Xmdls_inv_8 SS mdls_inv_6/IN mdls_inv_8/IN DD SS mdls_inv
Xring_100mV_buffer_0 ring_100mV_buffer_0/OUT mdls_inv_3/OUT DD SS ring_100mV_buffer
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_4HNDKD a_n500_n188# a_n660_n274# a_500_n100# a_n558_n100#
X0 a_500_n100# a_n500_n188# a_n558_n100# a_n660_n274# sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=5
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_C9VRMX a_n158_n250# a_n100_n338# a_100_n250# VSUBS
X0 a_100_n250# a_n100_n338# a_n158_n250# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
.ends

.subckt iref_2nA_igenerator Ip2 Ip1 Vg VCTAT SS
Xsky130_fd_pr__nfet_01v8_lvt_4HNDKD_0 VCTAT SS SS li_5063_n2421# sky130_fd_pr__nfet_01v8_lvt_4HNDKD
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_0 Ip2 Vg SS SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_1 SS SS SS SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_3 Ip1 Vg li_5063_n2421# SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_4 Ip1 Vg li_5063_n2421# SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_6 Ip2 Vg SS SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_7 SS SS SS SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_NTRJ8S a_200_n250# w_n294_n350# a_n200_n347# a_n258_n250#
X0 a_200_n250# a_n200_n347# a_n258_n250# w_n294_n350# sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_WCVK8S a_n200_n147# a_n258_n50# a_200_n50# w_n294_n150#
X0 a_200_n50# a_n200_n147# a_n258_n50# w_n294_n150# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
.ends

.subckt iref_2nA_mirrors Iref Ip2 Ip1 Vg DD SS
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_7 li_395_966# DD Ip1 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_6 li_1196_964# DD Ip1 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_8 m1_373_2671# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_9 m1_373_2671# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_40 m1_792_538# DD m1_792_538# m1_9767_755# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_30 m1_373_2671# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_31 Ip2 DD m1_792_538# m1_373_2671# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_20 Iref DD m1_792_538# li_5100_2660# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_42 m1_9767_755# DD m1_9767_755# DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_41 m1_792_538# DD m1_792_538# m1_9767_755# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_WCVK8S_0 DD DD DD DD sky130_fd_pr__pfet_01v8_lvt_WCVK8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_10 li_5100_2660# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_21 li_452_n361# DD m1_792_538# li_4299_2662# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_32 Ip2 DD m1_792_538# m1_373_2671# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_43 m1_9767_755# DD m1_9767_755# DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_WCVK8S_1 DD DD DD DD sky130_fd_pr__pfet_01v8_lvt_WCVK8S
Xsky130_fd_pr__pfet_01v8_lvt_WCVK8S_2 DD DD DD DD sky130_fd_pr__pfet_01v8_lvt_WCVK8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_22 li_5100_2660# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_11 li_4299_2662# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_33 m1_373_2671# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_WCVK8S_3 DD DD DD DD sky130_fd_pr__pfet_01v8_lvt_WCVK8S
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_10 m1_792_538# li_452_n361# SS SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_23 li_4299_2662# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_34 Ip2 DD m1_792_538# m1_373_2671# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_12 Ip2 DD m1_792_538# m1_373_2671# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_WCVK8S_4 DD DD DD DD sky130_fd_pr__pfet_01v8_lvt_WCVK8S
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_11 li_452_n361# li_452_n361# SS SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_35 m1_373_2671# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_WCVK8S_5 DD DD DD DD sky130_fd_pr__pfet_01v8_lvt_WCVK8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_13 Ip2 DD m1_792_538# m1_373_2671# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_12 li_452_n361# li_452_n361# SS SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_36 m1_373_2671# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_WCVK8S_6 DD DD DD DD sky130_fd_pr__pfet_01v8_lvt_WCVK8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_14 Iref DD m1_792_538# li_5100_2660# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_13 m1_792_538# li_452_n361# SS SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__pfet_01v8_lvt_WCVK8S_7 DD DD DD DD sky130_fd_pr__pfet_01v8_lvt_WCVK8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_37 Ip2 DD m1_792_538# m1_373_2671# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_26 Ip2 DD m1_792_538# m1_373_2671# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_15 li_452_n361# DD m1_792_538# li_4299_2662# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_14 Vg li_452_n361# SS SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_27 m1_373_2671# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_16 m1_373_2671# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_38 Ip2 DD m1_792_538# m1_373_2671# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_15 SS SS SS SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_39 m1_373_2671# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_18 Ip2 DD m1_792_538# m1_373_2671# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_17 Ip2 DD m1_792_538# m1_373_2671# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_8 SS SS SS SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_19 m1_373_2671# DD Ip2 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__nfet_01v8_lvt_C9VRMX_9 Vg li_452_n361# SS SS sky130_fd_pr__nfet_01v8_lvt_C9VRMX
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_0 Ip1 DD m1_792_538# li_395_966# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_1 Vg DD m1_792_538# li_1196_964# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_2 Vg DD m1_792_538# li_1196_964# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_3 Ip1 DD m1_792_538# li_395_966# sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_4 li_395_966# DD Ip1 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
Xsky130_fd_pr__pfet_01v8_lvt_NTRJ8S_5 li_1196_964# DD Ip1 DD sky130_fd_pr__pfet_01v8_lvt_NTRJ8S
.ends

.subckt iref_2nA_vref SS VREF DD
X0 VREF SS SS VREF sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X1 DD a_n1179_n2108# w_297_n2846# DD sky130_fd_pr__pfet_01v8 ad=0.687 pd=5.32 as=0.687 ps=5.32 w=2.37 l=4.38
X2 VREF SS SS VREF sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X3 DD DD a_n1179_n2108# DD sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X4 a_n1179_n2108# w_297_n2846# VREF DD sky130_fd_pr__pfet_01v8_lvt ad=0.995 pd=7.44 as=0.995 ps=7.44 w=3.43 l=2.77
X5 VREF SS SS VREF sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X6 w_297_n2846# w_297_n2846# SS w_297_n2846# sky130_fd_pr__pfet_01v8_lvt ad=0.255 pd=2.34 as=0.255 ps=2.34 w=0.88 l=6.97
X7 VREF SS SS VREF sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt iref_2nA DD IREF SS
Xiref_2nA_igenerator_0 iref_2nA_mirrors_0/Ip2 iref_2nA_mirrors_0/Ip1 iref_2nA_mirrors_0/Vg
+ iref_2nA_vref_0/VREF SS iref_2nA_igenerator
Xiref_2nA_mirrors_0 IREF iref_2nA_mirrors_0/Ip2 iref_2nA_mirrors_0/Ip1 iref_2nA_mirrors_0/Vg
+ DD SS iref_2nA_mirrors
Xiref_2nA_vref_0 SS iref_2nA_vref_0/VREF DD iref_2nA_vref
.ends

.subckt vref01 VREF DD SS
X0 SS a_n354_1346# VREF SS sky130_fd_pr__nfet_01v8 ad=0.238 pd=2.22 as=0.238 ps=2.22 w=0.82 l=1.05
X1 DD a_n354_1346# a_n354_1346# SS sky130_fd_pr__nfet_01v8_lvt ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.89
X2 VREF a_n354_1346# a_n354_1346# SS sky130_fd_pr__nfet_01v8_lvt ad=0.499 pd=4.02 as=0.499 ps=4.02 w=1.72 l=3.1
X3 VREF VREF VREF DD sky130_fd_pr__pfet_01v8_lvt ad=17.2 pd=38.4 as=8.6 ps=19.2 w=8.6 l=0.35
X4 DD a_n354_1346# a_n354_1346# SS sky130_fd_pr__nfet_01v8_lvt ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.89
.ends

.subckt pmu_circuits ldo_iref ldo_vs ring_out iref dd_02 dd_01 ldo_vb ldo_out vref
+ ss
Xldo_0 ldo_iref ss ldo_vb ldo_vs ldo_out dd_01 ldo
Xring_100mV_0 ss dd_02 ring_out ring_100mV
Xiref_2nA_0 dd_01 iref ss iref_2nA
Xvref01_0 vref dd_01 ss vref01
.ends

.subckt user_analog_proj_example pmu_circuits_0/iref pmu_circuits_0/dd_02 pmu_circuits_0/dd_01
+ pmu_circuits_0/ldo_vb pmu_circuits_0/ldo_iref pmu_circuits_0/ring_out pmu_circuits_0/ldo_vs
+ pmu_circuits_0/ldo_out VSUBS pmu_circuits_0/vref
Xpmu_circuits_0 pmu_circuits_0/ldo_iref pmu_circuits_0/ldo_vs pmu_circuits_0/ring_out
+ pmu_circuits_0/iref pmu_circuits_0/dd_02 pmu_circuits_0/dd_01 pmu_circuits_0/ldo_vb
+ pmu_circuits_0/ldo_out pmu_circuits_0/vref VSUBS pmu_circuits
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xuser_analog_proj_example_0 io_out[11] vdda1 vccd1 io_out[12] gpio_analog[7] gpio_analog[3]
+ io_out[16] io_out[15] vssa1 io_out[11] user_analog_proj_example
R0 io_oeb[15] vssd1 sky130_fd_pr__res_generic_m3 w=0.56 l=0.6
R1 io_analog[4] io_clamp_high[0] sky130_fd_pr__res_generic_m3 w=11 l=0.25
R2 vssd1 io_oeb[11] sky130_fd_pr__res_generic_m3 w=0.56 l=0.58
R3 vssa1 io_clamp_low[1] sky130_fd_pr__res_generic_m3 w=11 l=0.25
R4 io_oeb[16] vssd1 sky130_fd_pr__res_generic_m3 w=0.56 l=0.31
R5 vssa1 io_clamp_low[0] sky130_fd_pr__res_generic_m3 w=11 l=0.25
R6 vssd1 io_oeb[12] sky130_fd_pr__res_generic_m3 w=0.56 l=0.49
R7 vssa1 io_clamp_high[2] sky130_fd_pr__res_generic_m3 w=11 l=0.25
R8 vssa1 io_clamp_high[1] sky130_fd_pr__res_generic_m3 w=11 l=0.25
R9 vssa1 io_clamp_low[2] sky130_fd_pr__res_generic_m3 w=11 l=0.25
.ends


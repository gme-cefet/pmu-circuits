magic
tech sky130A
magscale 1 2
timestamp 1698329069
<< nwell >>
rect -1790 197 -945 2350
<< nmos >>
rect 916 864 1126 1028
<< pmoslvt >>
rect -1403 409 -1333 2129
<< nmoslvt >>
rect -266 1716 934 1894
rect -266 1346 934 1524
rect 28 756 648 1100
<< ndiff >>
rect -266 1940 934 1952
rect -266 1906 -254 1940
rect 922 1906 934 1940
rect -266 1894 934 1906
rect -266 1704 934 1716
rect -266 1670 -254 1704
rect 922 1670 934 1704
rect -266 1658 934 1670
rect -266 1570 934 1582
rect -266 1536 -254 1570
rect 922 1536 934 1570
rect -266 1524 934 1536
rect -266 1334 934 1346
rect -266 1300 -254 1334
rect 922 1300 934 1334
rect -266 1288 934 1300
rect -30 1088 28 1100
rect -30 768 -18 1088
rect 16 768 28 1088
rect -30 756 28 768
rect 648 1088 706 1100
rect 648 768 660 1088
rect 694 768 706 1088
rect 858 1016 916 1028
rect 858 876 870 1016
rect 904 876 916 1016
rect 858 864 916 876
rect 1126 1016 1184 1028
rect 1126 876 1138 1016
rect 1172 876 1184 1016
rect 1126 864 1184 876
rect 648 756 706 768
<< pdiff >>
rect -1603 2117 -1403 2129
rect -1603 421 -1449 2117
rect -1415 421 -1403 2117
rect -1603 409 -1403 421
rect -1333 2117 -1133 2129
rect -1333 421 -1321 2117
rect -1287 421 -1133 2117
rect -1333 409 -1133 421
<< ndiffc >>
rect -254 1906 922 1940
rect -254 1670 922 1704
rect -254 1536 922 1570
rect -254 1300 922 1334
rect -18 768 16 1088
rect 660 768 694 1088
rect 870 876 904 1016
rect 1138 876 1172 1016
<< pdiffc >>
rect -1449 421 -1415 2117
rect -1321 421 -1287 2117
<< psubdiff >>
rect -2152 2658 1826 2666
rect -2152 2642 -1860 2658
rect -1974 2501 -1860 2642
rect 1537 2642 1826 2658
rect 1537 2501 1648 2642
rect -696 2062 -576 2102
rect -622 2034 -576 2062
rect 1238 2062 1392 2102
rect 1238 2034 1318 2062
rect -622 496 -550 536
rect -696 468 -550 496
rect 1144 468 1220 536
rect 1264 496 1318 536
rect 1264 468 1392 496
rect -1974 41 1648 49
rect -1974 -83 -1870 41
rect -2152 -116 -1870 -83
rect 1527 -83 1648 41
rect 1527 -116 1826 -83
<< nsubdiff >>
rect -1754 2280 -1694 2314
rect -1041 2280 -981 2314
rect -1754 2254 -1720 2280
rect -1015 2254 -981 2280
rect -1754 267 -1720 293
rect -1015 267 -981 293
rect -1754 233 -1694 267
rect -1041 233 -981 267
<< psubdiffcont >>
rect -2152 -83 -1974 2642
rect -1860 2501 1537 2658
rect -696 496 -622 2062
rect -576 2034 1238 2102
rect -550 468 1144 536
rect 1220 468 1264 536
rect 1318 496 1392 2062
rect -1870 -116 1527 41
rect 1648 -83 1826 2642
<< nsubdiffcont >>
rect -1694 2280 -1041 2314
rect -1754 293 -1720 2254
rect -1015 293 -981 2254
rect -1694 233 -1041 267
<< poly >>
rect -1403 2210 -1333 2226
rect -1403 2176 -1387 2210
rect -1349 2176 -1333 2210
rect -1403 2129 -1333 2176
rect -1403 362 -1333 409
rect -1403 328 -1387 362
rect -1349 328 -1333 362
rect -1403 312 -1333 328
rect -354 1878 -266 1894
rect -354 1732 -338 1878
rect -304 1732 -266 1878
rect -354 1716 -266 1732
rect 934 1878 1022 1894
rect 934 1732 972 1878
rect 1006 1732 1022 1878
rect 934 1716 1022 1732
rect -354 1508 -266 1524
rect -354 1362 -338 1508
rect -304 1362 -266 1508
rect -354 1346 -266 1362
rect 934 1508 1022 1524
rect 934 1362 972 1508
rect 1006 1362 1022 1508
rect 934 1346 1022 1362
rect 28 1172 648 1188
rect 28 1138 44 1172
rect 632 1138 648 1172
rect 28 1100 648 1138
rect 916 1100 1126 1116
rect 916 1066 932 1100
rect 1110 1066 1126 1100
rect 916 1028 1126 1066
rect 916 826 1126 864
rect 916 792 932 826
rect 1110 792 1126 826
rect 916 776 1126 792
rect 28 718 648 756
rect 28 684 44 718
rect 632 684 648 718
rect 28 668 648 684
<< polycont >>
rect -1387 2176 -1349 2210
rect -1387 328 -1349 362
rect -338 1732 -304 1878
rect 972 1732 1006 1878
rect -338 1362 -304 1508
rect 972 1362 1006 1508
rect 44 1138 632 1172
rect 932 1066 1110 1100
rect 932 792 1110 826
rect 44 684 632 718
<< locali >>
rect -2152 2658 1826 2666
rect -2152 2642 -1860 2658
rect -1974 2501 -1860 2642
rect 1537 2642 1826 2658
rect 1537 2501 1648 2642
rect -1754 2280 -1694 2314
rect -1041 2280 -981 2314
rect -1754 2254 -1720 2280
rect -1015 2254 -981 2280
rect -1449 2176 -1387 2210
rect -1349 2176 -1287 2210
rect -1449 2117 -1415 2176
rect -1449 362 -1415 421
rect -1321 2117 -1287 2176
rect -1321 362 -1287 421
rect -1449 328 -1387 362
rect -1349 328 -1287 362
rect -1754 267 -1720 293
rect -696 2062 -576 2102
rect -981 1998 -840 2024
rect -981 1830 -970 1998
rect -869 1830 -840 1998
rect -981 1806 -840 1830
rect -622 2034 -576 2062
rect 1238 2062 1392 2102
rect 1238 2034 1318 2062
rect -270 1906 -254 1940
rect 922 1906 938 1940
rect -338 1878 -304 1894
rect -338 1716 -304 1732
rect 972 1878 1006 1894
rect 972 1716 1006 1732
rect -270 1670 -254 1704
rect 922 1670 938 1704
rect -270 1536 -254 1570
rect 922 1536 938 1570
rect -338 1508 -304 1524
rect -338 1346 -304 1362
rect 972 1508 1006 1524
rect 972 1346 1006 1362
rect -270 1300 -254 1334
rect 922 1300 938 1334
rect 28 1138 44 1172
rect 632 1138 648 1172
rect -18 1088 16 1104
rect -18 752 16 768
rect 660 1088 694 1104
rect 916 1066 932 1100
rect 1110 1066 1126 1100
rect 870 1016 904 1032
rect 870 860 904 876
rect 1138 1016 1318 1032
rect 1172 876 1318 1016
rect 1138 860 1318 876
rect 916 792 932 826
rect 1110 792 1126 826
rect 660 752 694 768
rect 28 684 44 718
rect 632 684 648 718
rect -622 496 -550 536
rect -696 468 -550 496
rect 1144 468 1220 536
rect 1264 496 1318 536
rect 1264 468 1392 496
rect -1015 267 -981 293
rect -1754 233 -1694 267
rect -1041 233 -981 267
rect -143 49 764 468
rect -1974 41 1648 49
rect -1974 -83 -1870 41
rect -2152 -116 -1870 -83
rect 1527 -83 1648 41
rect 1527 -116 1826 -83
<< viali >>
rect -1387 2176 -1349 2210
rect -1449 421 -1415 2117
rect -1321 421 -1287 2117
rect -1387 328 -1349 362
rect -970 1830 -869 1998
rect -254 1906 922 1940
rect -338 1732 -304 1878
rect 972 1732 1006 1878
rect -254 1670 922 1704
rect -254 1536 922 1570
rect -338 1362 -304 1508
rect 972 1362 1006 1508
rect -254 1300 922 1334
rect 44 1138 632 1172
rect -18 768 16 1088
rect 660 768 694 1088
rect 932 1066 1110 1100
rect 870 876 904 1016
rect 1138 876 1172 1016
rect 932 792 1110 826
rect 44 684 632 718
<< metal1 >>
rect -1449 2210 -1287 2226
rect -1449 2176 -1387 2210
rect -1349 2176 -1287 2210
rect -1399 2170 -1337 2176
rect -1455 2117 -1409 2129
rect -1455 421 -1449 2117
rect -1415 421 -1409 2117
rect -1455 409 -1409 421
rect -1327 2117 -1281 2129
rect -1327 421 -1321 2117
rect -1287 825 -1281 2117
rect -999 1998 4 2024
rect -999 1830 -970 1998
rect -869 1986 4 1998
rect -869 1830 -706 1986
rect -999 1806 -706 1830
rect -590 1946 4 1986
rect -590 1944 934 1946
rect -590 1618 -444 1944
rect -266 1940 934 1944
rect -266 1906 -254 1940
rect 922 1906 934 1940
rect -266 1900 934 1906
rect -400 1878 -298 1890
rect -400 1732 -390 1878
rect -304 1732 -298 1878
rect -400 1720 -298 1732
rect 966 1878 1156 1890
rect 966 1732 972 1878
rect 1058 1732 1156 1878
rect 966 1720 1156 1732
rect -266 1704 934 1710
rect -266 1670 -254 1704
rect 922 1670 934 1704
rect -266 1664 934 1670
rect 878 1658 934 1664
rect 1068 1658 1086 1720
rect 878 1622 1086 1658
rect -590 1576 4 1618
rect -266 1570 934 1576
rect -266 1536 -254 1570
rect 922 1536 934 1570
rect -266 1530 934 1536
rect 1068 1522 1086 1622
rect 1142 1522 1156 1720
rect 1068 1520 1156 1522
rect -400 1508 -298 1520
rect -400 1362 -390 1508
rect -304 1362 -298 1508
rect -400 1350 -298 1362
rect 966 1508 1156 1520
rect 966 1362 972 1508
rect 1058 1362 1156 1508
rect 966 1350 1156 1362
rect -400 1224 -358 1350
rect -266 1334 934 1340
rect -266 1300 -254 1334
rect 922 1300 934 1334
rect -266 1294 934 1300
rect -266 1224 -158 1294
rect -400 1176 -158 1224
rect -266 1014 -158 1176
rect 32 1248 644 1294
rect 1080 1248 1156 1350
rect 32 1198 1156 1248
rect 32 1172 644 1198
rect 32 1138 44 1172
rect 632 1138 644 1172
rect 32 1132 644 1138
rect 920 1100 1156 1198
rect -24 1088 22 1100
rect -24 1014 -18 1088
rect -266 850 -18 1014
rect -734 825 -488 840
rect -1287 814 -488 825
rect -1287 752 -734 814
rect -534 752 -488 814
rect -1287 747 -488 752
rect -1287 421 -1281 747
rect -734 722 -488 747
rect -266 678 -136 850
rect -24 768 -18 850
rect 16 768 22 1088
rect -24 756 22 768
rect 654 1088 700 1100
rect 654 768 660 1088
rect 694 1028 700 1088
rect 920 1066 932 1100
rect 1110 1066 1156 1100
rect 920 1060 1156 1066
rect 694 1016 910 1028
rect 694 1006 870 1016
rect 694 882 730 1006
rect 832 882 870 1006
rect 694 876 870 882
rect 904 876 910 1016
rect 694 864 910 876
rect 1132 1016 1178 1028
rect 1132 876 1138 1016
rect 1172 876 1178 1016
rect 1132 864 1178 876
rect 694 768 700 864
rect 654 756 700 768
rect 920 826 1122 832
rect 920 792 932 826
rect 1110 792 1122 826
rect 32 718 644 724
rect 32 684 44 718
rect 632 684 644 718
rect 32 678 644 684
rect 920 678 1122 792
rect -266 620 1122 678
rect -1327 409 -1281 421
rect -1449 362 -1287 368
rect -1449 328 -1387 362
rect -1349 328 -1287 362
rect -1449 322 -1287 328
<< via1 >>
rect -390 1732 -338 1878
rect 1006 1732 1058 1878
rect 1086 1522 1142 1720
rect -390 1362 -338 1508
rect 1006 1362 1058 1508
rect -734 752 -534 814
rect 730 882 832 1006
<< metal2 >>
rect -400 1878 -298 1890
rect -400 1732 -390 1878
rect -338 1732 -298 1878
rect -400 1720 -298 1732
rect 966 1878 1156 1890
rect 966 1732 1006 1878
rect 1058 1732 1156 1878
rect 966 1720 1156 1732
rect -400 1520 -344 1720
rect 1012 1522 1086 1720
rect 1142 1522 1156 1720
rect 1012 1520 1156 1522
rect -400 1508 -298 1520
rect -400 1362 -390 1508
rect -338 1362 -298 1508
rect -400 1350 -298 1362
rect 966 1508 1156 1520
rect 966 1362 1006 1508
rect 1058 1362 1156 1508
rect 966 1350 1156 1362
rect 706 1006 858 1028
rect 706 882 730 1006
rect 832 882 858 1006
rect 706 864 858 882
rect -734 814 -446 840
rect -534 752 -446 814
rect -734 722 -446 752
rect -504 628 -446 722
rect 756 628 858 864
rect -504 558 858 628
<< labels >>
flabel metal2 -484 566 -416 614 0 FreeSans 1600 0 0 0 VREF
port 0 nsew
flabel metal1 -548 1916 -480 1964 0 FreeSans 1600 0 0 0 DD
port 1 nsew
flabel locali 1230 908 1298 956 0 FreeSans 1600 0 0 0 SS
port 2 nsew
<< end >>

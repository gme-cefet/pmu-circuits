magic
tech sky130A
magscale 1 2
timestamp 1697410379
use pmu_circuits  pmu_circuits_0
timestamp 1697410379
transform 1 0 11036 0 1 -3638
box -1074 5482 18938 20761
<< end >>

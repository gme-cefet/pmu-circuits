magic
tech sky130A
magscale 1 2
timestamp 1697410379
<< locali >>
rect -1047 19784 18654 20384
rect -1047 7299 -494 19784
rect 5507 19629 12606 19784
rect 16247 17627 17282 19784
rect 16247 17621 16975 17627
rect 11510 15672 11938 16174
rect -1047 7076 2091 7299
rect 5959 7076 12804 7245
rect 14590 7076 15868 7365
rect -1047 6476 18788 7076
rect -1047 6466 -494 6476
<< metal1 >>
rect 11103 17945 12417 17992
rect 11103 17720 11162 17945
rect 12344 17720 12417 17945
rect 11103 17676 12417 17720
rect 13052 16088 13638 20761
rect 12650 15851 13638 16088
rect 14338 18091 15837 18358
rect 14338 14470 14605 18091
rect 15570 17552 15837 18091
rect 15570 17460 15931 17552
rect 15798 17362 15931 17460
rect 13599 14255 14605 14470
rect 13597 13886 18539 14255
rect 4766 9676 5354 9772
rect 4766 7246 4854 9676
rect 5270 7246 5354 9676
rect 4766 7166 5354 7246
rect 4766 6140 5352 7166
rect 13599 6140 14090 13886
rect 17989 13735 18511 13886
rect 18067 10565 18686 10994
rect 18401 10009 18782 10214
rect 16311 7296 16465 7327
rect 16311 7117 18938 7296
rect -726 5482 18815 6140
<< via1 >>
rect 11162 17720 12344 17945
rect 4854 7246 5270 9676
<< metal2 >>
rect 12233 17992 12413 20748
rect 11103 17945 12417 17992
rect 11103 17720 11162 17945
rect 12344 17720 12417 17945
rect 11103 17676 12417 17720
rect 16482 15937 16626 16160
rect 16482 15844 18576 15937
rect 16483 15706 18576 15844
rect 4766 9676 5354 9760
rect 4766 7781 4854 9676
rect 4456 7246 4854 7781
rect 5270 7246 5354 9676
rect 4456 7243 5354 7246
rect 4766 7166 5354 7243
<< metal3 >>
rect -1074 8423 461 9174
rect 18391 8894 18870 9125
use iref_2nA  iref_2nA_0
timestamp 1697064583
transform 0 1 4468 -1 0 16274
box -3409 -5056 9048 205
use ldo  ldo_0
timestamp 1697396974
transform 1 0 5724 0 1 17576
box 8574 -10258 12913 -3712
use ring_100mV  ring_100mV_0
timestamp 1697065484
transform 1 0 4604 0 1 12805
box 848 -5593 8961 6935
use vref01  vref01_0
timestamp 1697409234
transform 1 0 16504 0 1 15556
box -1790 197 1392 2350
<< labels >>
flabel metal1 17837 5640 18206 5982 0 FreeSans 4800 0 0 0 dd_01
flabel metal2 12247 20563 12392 20714 0 FreeSans 4800 0 0 0 ring_out
flabel metal1 13288 17947 13433 18098 0 FreeSans 4800 90 0 0 dd_02
flabel metal2 18164 15752 18309 15903 0 FreeSans 4800 0 0 0 vref
flabel metal3 -956 8734 -811 8885 0 FreeSans 4800 0 0 0 iref
flabel metal1 18510 10716 18655 10867 0 FreeSans 4800 0 0 0 ldo_out
flabel metal1 18604 10029 18749 10180 0 FreeSans 4800 0 0 0 ldo_vs
flabel metal3 18678 8947 18823 9098 0 FreeSans 4800 0 0 0 ldo_vb
flabel metal1 18520 7171 18648 7255 0 FreeSans 4800 0 0 0 ldo_iref
flabel locali -728 6674 -273 7080 0 FreeSans 4800 0 0 0 ss
<< end >>

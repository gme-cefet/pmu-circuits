magic
tech sky130A
timestamp 1697035654
<< nmoslvt >>
rect -40 -275 40 275
<< ndiff >>
rect -69 269 -40 275
rect -69 -269 -63 269
rect -46 -269 -40 269
rect -69 -275 -40 -269
rect 40 269 69 275
rect 40 -269 46 269
rect 63 -269 69 269
rect 40 -275 69 -269
<< ndiffc >>
rect -63 -269 -46 269
rect 46 -269 63 269
<< poly >>
rect -40 311 40 319
rect -40 294 -32 311
rect 32 294 40 311
rect -40 275 40 294
rect -40 -294 40 -275
rect -40 -311 -32 -294
rect 32 -311 40 -294
rect -40 -319 40 -311
<< polycont >>
rect -32 294 32 311
rect -32 -311 32 -294
<< locali >>
rect -40 294 -32 311
rect 32 294 40 311
rect -63 269 -46 277
rect -63 -277 -46 -269
rect 46 269 63 277
rect 46 -277 63 -269
rect -40 -311 -32 -294
rect 32 -311 40 -294
<< viali >>
rect -32 294 32 311
rect -63 -269 -46 269
rect 46 -269 63 269
rect -32 -311 32 -294
<< metal1 >>
rect -38 311 38 314
rect -38 294 -32 311
rect 32 294 38 311
rect -38 291 38 294
rect -66 269 -43 275
rect -66 -269 -63 269
rect -46 -269 -43 269
rect -66 -275 -43 -269
rect 43 269 66 275
rect 43 -269 46 269
rect 63 -269 66 269
rect 43 -275 66 -269
rect -38 -294 38 -291
rect -38 -311 -32 -294
rect 32 -311 38 -294
rect -38 -314 38 -311
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.5 l 0.8 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

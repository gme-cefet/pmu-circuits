magic
tech sky130A
magscale 1 2
timestamp 1698332589
<< nwell >>
rect 2727 19433 4410 19449
rect 1021 15357 4410 19433
rect 9044 16669 12374 17667
rect 14714 15753 15559 17906
rect -382 12384 2364 12876
rect 583 11504 2369 12118
rect 205 9873 2393 11240
rect 937 7748 2478 9461
rect 2847 9255 4410 15357
rect 937 7747 2469 7748
rect 2842 7542 4410 9255
rect 8825 7392 10192 15722
rect 14728 12421 17941 13714
rect 16867 11031 18339 11497
rect 16807 9133 18478 10477
<< pwell >>
rect 463 13319 1855 13939
rect 14352 9170 15030 11884
<< nmos >>
rect 17420 16420 17630 16584
<< pmos >>
rect -163 12580 237 12680
rect 473 12580 873 12680
rect 1109 12580 1509 12680
rect 1745 12580 2145 12680
rect 1321 10125 2197 10599
rect 14982 12678 15160 13456
rect 15482 12678 15660 13456
rect 15982 12678 16160 13456
rect 16482 12678 16660 13456
rect 16982 12678 17160 13456
rect 17482 12678 17660 13456
<< pmoslvt >>
rect 1386 19098 1786 19198
rect 2086 19098 2486 19198
rect 1386 18314 1786 18814
rect 2086 18314 2486 18814
rect 1386 17530 1786 18030
rect 2086 17530 2486 18030
rect 1386 16746 1786 17246
rect 2086 16746 2486 17246
rect 1386 15962 1786 16462
rect 2086 15962 2486 16462
rect 1386 15578 1786 15678
rect 2086 15578 2486 15678
rect 779 11723 2173 11899
rect 401 10311 955 10997
rect 1395 10891 2195 10991
rect 1155 8752 1555 9252
rect 1855 8752 2255 9252
rect 1155 7968 1555 8468
rect 1855 7968 2255 8468
rect 3082 19114 3482 19214
rect 3782 19114 4182 19214
rect 3082 18330 3482 18830
rect 3782 18330 4182 18830
rect 3082 17546 3482 18046
rect 3782 17546 4182 18046
rect 3082 16762 3482 17262
rect 3782 16762 4182 17262
rect 3082 15978 3482 16478
rect 3782 15978 4182 16478
rect 3082 15194 3482 15694
rect 3782 15194 4182 15694
rect 3082 14410 3482 14910
rect 3782 14410 4182 14910
rect 3082 13626 3482 14126
rect 3782 13626 4182 14126
rect 3082 12842 3482 13342
rect 3782 12842 4182 13342
rect 3082 12058 3482 12558
rect 3782 12058 4182 12558
rect 3082 11274 3482 11774
rect 3782 11274 4182 11774
rect 3082 10490 3482 10990
rect 3782 10490 4182 10990
rect 3082 9706 3482 10206
rect 3782 9706 4182 10206
rect 3082 8922 3482 9422
rect 3782 8922 4182 9422
rect 3082 8138 3482 8638
rect 3782 8138 4182 8638
rect 3082 7754 3482 7854
rect 3782 7754 4182 7854
rect 9414 17114 9574 17314
rect 9814 17114 9974 17314
rect 10673 17085 10833 17285
rect 11073 17085 11233 17285
rect 11473 17085 11633 17285
rect 11873 17085 12033 17285
rect 9063 15346 9263 15506
rect 9063 14938 9263 15098
rect 9063 14252 9263 14652
rect 9754 15346 9954 15506
rect 9754 14938 9954 15098
rect 9754 14252 9954 14652
rect 9063 13680 9263 13840
rect 9063 13272 9263 13432
rect 9063 12586 9263 12986
rect 9754 13680 9954 13840
rect 9754 13272 9954 13432
rect 9754 12586 9954 12986
rect 9063 12014 9263 12174
rect 9063 11606 9263 11766
rect 9063 10920 9263 11320
rect 9754 12014 9954 12174
rect 9754 11606 9954 11766
rect 9754 10920 9954 11320
rect 9063 10348 9263 10508
rect 9063 9940 9263 10100
rect 9063 9254 9263 9654
rect 9754 10348 9954 10508
rect 9754 9940 9954 10100
rect 9754 9254 9954 9654
rect 9063 8682 9263 8842
rect 9063 8274 9263 8434
rect 9063 7588 9263 7988
rect 9754 8682 9954 8842
rect 9754 8274 9954 8434
rect 9754 7588 9954 7988
rect 15101 15965 15171 17685
rect 17086 11227 18120 11301
rect 17029 9980 18243 10234
rect 17029 9380 18243 9634
<< nmoslvt >>
rect -81 18783 419 18983
rect -81 18367 419 18567
rect -81 17951 419 18151
rect -81 17535 419 17735
rect -81 17119 419 17319
rect -81 16703 419 16903
rect -81 16287 419 16487
rect -81 15871 419 16071
rect 54 14113 254 14613
rect 470 14113 670 14613
rect 886 14113 1086 14613
rect 1302 14113 1502 14613
rect 1718 14113 1918 14613
rect 2134 14113 2334 14613
rect 659 13529 1659 13729
rect 5891 18167 6051 19267
rect 6291 18167 6451 19267
rect 6691 18167 6851 19267
rect 7091 18167 7251 19267
rect 7491 18167 7651 19267
rect 7891 18167 8051 19267
rect 8291 18167 8451 19267
rect 8691 18167 8851 19267
rect 9091 18167 9251 19267
rect 9491 18167 9651 19267
rect 9891 18167 10051 19267
rect 10291 18167 10451 19267
rect 10691 18167 10851 19267
rect 11091 18167 11251 19267
rect 11491 18167 11651 19267
rect 11891 18167 12051 19267
rect 5770 16467 5930 17567
rect 6170 16467 6330 17567
rect 6570 16467 6730 17567
rect 6970 16467 7130 17567
rect 7370 16467 7530 17567
rect 7770 16467 7930 17567
rect 8170 16467 8330 17567
rect 8570 16467 8730 17567
rect 5930 15315 7030 15475
rect 7406 15351 8506 15431
rect 5930 14955 7030 15115
rect 7406 15053 8506 15133
rect 5930 14595 7030 14755
rect 7376 14651 8476 14851
rect 5930 14235 7030 14395
rect 7376 14227 8476 14427
rect 10511 15351 11611 15431
rect 11987 15315 13087 15475
rect 10511 15053 11611 15133
rect 11987 14955 13087 15115
rect 10541 14651 11641 14851
rect 11987 14595 13087 14755
rect 10541 14227 11641 14427
rect 11987 14235 13087 14395
rect 5930 13649 7030 13809
rect 7406 13685 8506 13765
rect 5930 13289 7030 13449
rect 7406 13387 8506 13467
rect 5930 12929 7030 13089
rect 7376 12985 8476 13185
rect 5930 12569 7030 12729
rect 7376 12561 8476 12761
rect 10511 13685 11611 13765
rect 11987 13649 13087 13809
rect 10511 13387 11611 13467
rect 11987 13289 13087 13449
rect 10541 12985 11641 13185
rect 11987 12929 13087 13089
rect 10541 12561 11641 12761
rect 11987 12569 13087 12729
rect 5930 11983 7030 12143
rect 7406 12019 8506 12099
rect 5930 11623 7030 11783
rect 7406 11721 8506 11801
rect 5930 11263 7030 11423
rect 7376 11319 8476 11519
rect 5930 10903 7030 11063
rect 7376 10895 8476 11095
rect 10511 12019 11611 12099
rect 11987 11983 13087 12143
rect 10511 11721 11611 11801
rect 11987 11623 13087 11783
rect 10541 11319 11641 11519
rect 11987 11263 13087 11423
rect 10541 10895 11641 11095
rect 11987 10903 13087 11063
rect 5930 10317 7030 10477
rect 7406 10353 8506 10433
rect 5930 9957 7030 10117
rect 7406 10055 8506 10135
rect 5930 9597 7030 9757
rect 7376 9653 8476 9853
rect 5930 9237 7030 9397
rect 7376 9229 8476 9429
rect 10511 10353 11611 10433
rect 11987 10317 13087 10477
rect 10511 10055 11611 10135
rect 11987 9957 13087 10117
rect 10541 9653 11641 9853
rect 11987 9597 13087 9757
rect 10541 9229 11641 9429
rect 11987 9237 13087 9397
rect 5930 8651 7030 8811
rect 7406 8687 8506 8767
rect 5930 8291 7030 8451
rect 7406 8389 8506 8469
rect 5930 7931 7030 8091
rect 7376 7987 8476 8187
rect 5930 7571 7030 7731
rect 7376 7563 8476 7763
rect 10511 8687 11611 8767
rect 11987 8651 13087 8811
rect 10511 8389 11611 8469
rect 11987 8291 13087 8451
rect 10541 7987 11641 8187
rect 11987 7931 13087 8091
rect 10541 7563 11641 7763
rect 11987 7571 13087 7731
rect 16238 17272 17438 17450
rect 16238 16902 17438 17080
rect 16532 16312 17152 16656
rect 14548 10636 14834 11674
rect 14548 9380 14834 10418
rect 14522 7578 14654 8598
rect 14922 7578 15054 8598
rect 15322 7578 15454 8598
rect 15722 7578 15854 8598
rect 16122 7578 16254 8598
rect 16522 7578 16654 8598
rect 16922 7578 17054 8598
rect 17322 7578 17454 8598
rect 17722 7578 17854 8598
rect 18122 7578 18254 8598
<< ndiff >>
rect -81 19029 419 19041
rect -81 18995 -69 19029
rect 407 18995 419 19029
rect -81 18983 419 18995
rect -81 18771 419 18783
rect -81 18737 -69 18771
rect 407 18737 419 18771
rect -81 18725 419 18737
rect -81 18613 419 18625
rect -81 18579 -69 18613
rect 407 18579 419 18613
rect -81 18567 419 18579
rect -81 18355 419 18367
rect -81 18321 -69 18355
rect 407 18321 419 18355
rect -81 18309 419 18321
rect -81 18197 419 18209
rect -81 18163 -69 18197
rect 407 18163 419 18197
rect -81 18151 419 18163
rect -81 17939 419 17951
rect -81 17905 -69 17939
rect 407 17905 419 17939
rect -81 17893 419 17905
rect -81 17781 419 17793
rect -81 17747 -69 17781
rect 407 17747 419 17781
rect -81 17735 419 17747
rect -81 17523 419 17535
rect -81 17489 -69 17523
rect 407 17489 419 17523
rect -81 17477 419 17489
rect -81 17365 419 17377
rect -81 17331 -69 17365
rect 407 17331 419 17365
rect -81 17319 419 17331
rect -81 17107 419 17119
rect -81 17073 -69 17107
rect 407 17073 419 17107
rect -81 17061 419 17073
rect -81 16949 419 16961
rect -81 16915 -69 16949
rect 407 16915 419 16949
rect -81 16903 419 16915
rect -81 16691 419 16703
rect -81 16657 -69 16691
rect 407 16657 419 16691
rect -81 16645 419 16657
rect -81 16533 419 16545
rect -81 16499 -69 16533
rect 407 16499 419 16533
rect -81 16487 419 16499
rect -81 16275 419 16287
rect -81 16241 -69 16275
rect 407 16241 419 16275
rect -81 16229 419 16241
rect -81 16117 419 16129
rect -81 16083 -69 16117
rect 407 16083 419 16117
rect -81 16071 419 16083
rect -81 15859 419 15871
rect -81 15825 -69 15859
rect 407 15825 419 15859
rect -81 15813 419 15825
rect -4 14601 54 14613
rect -4 14125 8 14601
rect 42 14125 54 14601
rect -4 14113 54 14125
rect 254 14601 312 14613
rect 254 14125 266 14601
rect 300 14125 312 14601
rect 254 14113 312 14125
rect 412 14601 470 14613
rect 412 14125 424 14601
rect 458 14125 470 14601
rect 412 14113 470 14125
rect 670 14601 728 14613
rect 670 14125 682 14601
rect 716 14125 728 14601
rect 670 14113 728 14125
rect 828 14601 886 14613
rect 828 14125 840 14601
rect 874 14125 886 14601
rect 828 14113 886 14125
rect 1086 14601 1144 14613
rect 1086 14125 1098 14601
rect 1132 14125 1144 14601
rect 1086 14113 1144 14125
rect 1244 14601 1302 14613
rect 1244 14125 1256 14601
rect 1290 14125 1302 14601
rect 1244 14113 1302 14125
rect 1502 14601 1560 14613
rect 1502 14125 1514 14601
rect 1548 14125 1560 14601
rect 1502 14113 1560 14125
rect 1660 14601 1718 14613
rect 1660 14125 1672 14601
rect 1706 14125 1718 14601
rect 1660 14113 1718 14125
rect 1918 14601 1976 14613
rect 1918 14125 1930 14601
rect 1964 14125 1976 14601
rect 1918 14113 1976 14125
rect 2076 14601 2134 14613
rect 2076 14125 2088 14601
rect 2122 14125 2134 14601
rect 2076 14113 2134 14125
rect 2334 14601 2392 14613
rect 2334 14125 2346 14601
rect 2380 14125 2392 14601
rect 2334 14113 2392 14125
rect 601 13717 659 13729
rect 601 13541 613 13717
rect 647 13541 659 13717
rect 601 13529 659 13541
rect 1659 13717 1717 13729
rect 1659 13541 1671 13717
rect 1705 13541 1717 13717
rect 1659 13529 1717 13541
rect 5833 19255 5891 19267
rect 5833 18179 5845 19255
rect 5879 18179 5891 19255
rect 5833 18167 5891 18179
rect 6051 19255 6109 19267
rect 6051 18179 6063 19255
rect 6097 18179 6109 19255
rect 6051 18167 6109 18179
rect 6233 19255 6291 19267
rect 6233 18179 6245 19255
rect 6279 18179 6291 19255
rect 6233 18167 6291 18179
rect 6451 19255 6509 19267
rect 6451 18179 6463 19255
rect 6497 18179 6509 19255
rect 6451 18167 6509 18179
rect 6633 19255 6691 19267
rect 6633 18179 6645 19255
rect 6679 18179 6691 19255
rect 6633 18167 6691 18179
rect 6851 19255 6909 19267
rect 6851 18179 6863 19255
rect 6897 18179 6909 19255
rect 6851 18167 6909 18179
rect 7033 19255 7091 19267
rect 7033 18179 7045 19255
rect 7079 18179 7091 19255
rect 7033 18167 7091 18179
rect 7251 19255 7309 19267
rect 7251 18179 7263 19255
rect 7297 18179 7309 19255
rect 7251 18167 7309 18179
rect 7433 19255 7491 19267
rect 7433 18179 7445 19255
rect 7479 18179 7491 19255
rect 7433 18167 7491 18179
rect 7651 19255 7709 19267
rect 7651 18179 7663 19255
rect 7697 18179 7709 19255
rect 7651 18167 7709 18179
rect 7833 19255 7891 19267
rect 7833 18179 7845 19255
rect 7879 18179 7891 19255
rect 7833 18167 7891 18179
rect 8051 19255 8109 19267
rect 8051 18179 8063 19255
rect 8097 18179 8109 19255
rect 8051 18167 8109 18179
rect 8233 19255 8291 19267
rect 8233 18179 8245 19255
rect 8279 18179 8291 19255
rect 8233 18167 8291 18179
rect 8451 19255 8509 19267
rect 8451 18179 8463 19255
rect 8497 18179 8509 19255
rect 8451 18167 8509 18179
rect 8633 19255 8691 19267
rect 8633 18179 8645 19255
rect 8679 18179 8691 19255
rect 8633 18167 8691 18179
rect 8851 19255 8909 19267
rect 8851 18179 8863 19255
rect 8897 18179 8909 19255
rect 8851 18167 8909 18179
rect 9033 19255 9091 19267
rect 9033 18179 9045 19255
rect 9079 18179 9091 19255
rect 9033 18167 9091 18179
rect 9251 19255 9309 19267
rect 9251 18179 9263 19255
rect 9297 18179 9309 19255
rect 9251 18167 9309 18179
rect 9433 19255 9491 19267
rect 9433 18179 9445 19255
rect 9479 18179 9491 19255
rect 9433 18167 9491 18179
rect 9651 19255 9709 19267
rect 9651 18179 9663 19255
rect 9697 18179 9709 19255
rect 9651 18167 9709 18179
rect 9833 19255 9891 19267
rect 9833 18179 9845 19255
rect 9879 18179 9891 19255
rect 9833 18167 9891 18179
rect 10051 19255 10109 19267
rect 10051 18179 10063 19255
rect 10097 18179 10109 19255
rect 10051 18167 10109 18179
rect 10233 19255 10291 19267
rect 10233 18179 10245 19255
rect 10279 18179 10291 19255
rect 10233 18167 10291 18179
rect 10451 19255 10509 19267
rect 10451 18179 10463 19255
rect 10497 18179 10509 19255
rect 10451 18167 10509 18179
rect 10633 19255 10691 19267
rect 10633 18179 10645 19255
rect 10679 18179 10691 19255
rect 10633 18167 10691 18179
rect 10851 19255 10909 19267
rect 10851 18179 10863 19255
rect 10897 18179 10909 19255
rect 10851 18167 10909 18179
rect 11033 19255 11091 19267
rect 11033 18179 11045 19255
rect 11079 18179 11091 19255
rect 11033 18167 11091 18179
rect 11251 19255 11309 19267
rect 11251 18179 11263 19255
rect 11297 18179 11309 19255
rect 11251 18167 11309 18179
rect 11433 19255 11491 19267
rect 11433 18179 11445 19255
rect 11479 18179 11491 19255
rect 11433 18167 11491 18179
rect 11651 19255 11709 19267
rect 11651 18179 11663 19255
rect 11697 18179 11709 19255
rect 11651 18167 11709 18179
rect 11833 19255 11891 19267
rect 11833 18179 11845 19255
rect 11879 18179 11891 19255
rect 11833 18167 11891 18179
rect 12051 19255 12109 19267
rect 12051 18179 12063 19255
rect 12097 18179 12109 19255
rect 12051 18167 12109 18179
rect 5712 17555 5770 17567
rect 5712 16479 5724 17555
rect 5758 16479 5770 17555
rect 5712 16467 5770 16479
rect 5930 17555 5988 17567
rect 5930 16479 5942 17555
rect 5976 16479 5988 17555
rect 5930 16467 5988 16479
rect 6112 17555 6170 17567
rect 6112 16479 6124 17555
rect 6158 16479 6170 17555
rect 6112 16467 6170 16479
rect 6330 17555 6388 17567
rect 6330 16479 6342 17555
rect 6376 16479 6388 17555
rect 6330 16467 6388 16479
rect 6512 17555 6570 17567
rect 6512 16479 6524 17555
rect 6558 16479 6570 17555
rect 6512 16467 6570 16479
rect 6730 17555 6788 17567
rect 6730 16479 6742 17555
rect 6776 16479 6788 17555
rect 6730 16467 6788 16479
rect 6912 17555 6970 17567
rect 6912 16479 6924 17555
rect 6958 16479 6970 17555
rect 6912 16467 6970 16479
rect 7130 17555 7188 17567
rect 7130 16479 7142 17555
rect 7176 16479 7188 17555
rect 7130 16467 7188 16479
rect 7312 17555 7370 17567
rect 7312 16479 7324 17555
rect 7358 16479 7370 17555
rect 7312 16467 7370 16479
rect 7530 17555 7588 17567
rect 7530 16479 7542 17555
rect 7576 16479 7588 17555
rect 7530 16467 7588 16479
rect 7712 17555 7770 17567
rect 7712 16479 7724 17555
rect 7758 16479 7770 17555
rect 7712 16467 7770 16479
rect 7930 17555 7988 17567
rect 7930 16479 7942 17555
rect 7976 16479 7988 17555
rect 7930 16467 7988 16479
rect 8112 17555 8170 17567
rect 8112 16479 8124 17555
rect 8158 16479 8170 17555
rect 8112 16467 8170 16479
rect 8330 17555 8388 17567
rect 8330 16479 8342 17555
rect 8376 16479 8388 17555
rect 8330 16467 8388 16479
rect 8512 17555 8570 17567
rect 8512 16479 8524 17555
rect 8558 16479 8570 17555
rect 8512 16467 8570 16479
rect 8730 17555 8788 17567
rect 8730 16479 8742 17555
rect 8776 16479 8788 17555
rect 8730 16467 8788 16479
rect 5930 15521 7030 15533
rect 5930 15487 5942 15521
rect 7018 15487 7030 15521
rect 5930 15475 7030 15487
rect 7406 15477 8506 15489
rect 7406 15443 7418 15477
rect 8494 15443 8506 15477
rect 7406 15431 8506 15443
rect 7406 15339 8506 15351
rect 5930 15303 7030 15315
rect 5930 15269 5942 15303
rect 7018 15269 7030 15303
rect 7406 15305 7418 15339
rect 8494 15305 8506 15339
rect 7406 15293 8506 15305
rect 5930 15257 7030 15269
rect 7406 15179 8506 15191
rect 5930 15161 7030 15173
rect 5930 15127 5942 15161
rect 7018 15127 7030 15161
rect 7406 15145 7418 15179
rect 8494 15145 8506 15179
rect 7406 15133 8506 15145
rect 5930 15115 7030 15127
rect 7406 15041 8506 15053
rect 7406 15007 7418 15041
rect 8494 15007 8506 15041
rect 7406 14995 8506 15007
rect 5930 14943 7030 14955
rect 5930 14909 5942 14943
rect 7018 14909 7030 14943
rect 5930 14897 7030 14909
rect 7376 14897 8476 14909
rect 7376 14863 7388 14897
rect 8464 14863 8476 14897
rect 7376 14851 8476 14863
rect 5930 14801 7030 14813
rect 5930 14767 5942 14801
rect 7018 14767 7030 14801
rect 5930 14755 7030 14767
rect 7376 14639 8476 14651
rect 7376 14605 7388 14639
rect 8464 14605 8476 14639
rect 5930 14583 7030 14595
rect 7376 14593 8476 14605
rect 5930 14549 5942 14583
rect 7018 14549 7030 14583
rect 5930 14537 7030 14549
rect 7376 14473 8476 14485
rect 5930 14441 7030 14453
rect 5930 14407 5942 14441
rect 7018 14407 7030 14441
rect 7376 14439 7388 14473
rect 8464 14439 8476 14473
rect 7376 14427 8476 14439
rect 5930 14395 7030 14407
rect 5930 14223 7030 14235
rect 5930 14189 5942 14223
rect 7018 14189 7030 14223
rect 5930 14177 7030 14189
rect 7376 14215 8476 14227
rect 7376 14181 7388 14215
rect 8464 14181 8476 14215
rect 7376 14169 8476 14181
rect 11987 15521 13087 15533
rect 10511 15477 11611 15489
rect 10511 15443 10523 15477
rect 11599 15443 11611 15477
rect 11987 15487 11999 15521
rect 13075 15487 13087 15521
rect 11987 15475 13087 15487
rect 10511 15431 11611 15443
rect 10511 15339 11611 15351
rect 10511 15305 10523 15339
rect 11599 15305 11611 15339
rect 10511 15293 11611 15305
rect 11987 15303 13087 15315
rect 11987 15269 11999 15303
rect 13075 15269 13087 15303
rect 11987 15257 13087 15269
rect 10511 15179 11611 15191
rect 10511 15145 10523 15179
rect 11599 15145 11611 15179
rect 10511 15133 11611 15145
rect 11987 15161 13087 15173
rect 11987 15127 11999 15161
rect 13075 15127 13087 15161
rect 11987 15115 13087 15127
rect 10511 15041 11611 15053
rect 10511 15007 10523 15041
rect 11599 15007 11611 15041
rect 10511 14995 11611 15007
rect 11987 14943 13087 14955
rect 11987 14909 11999 14943
rect 13075 14909 13087 14943
rect 10541 14897 11641 14909
rect 11987 14897 13087 14909
rect 10541 14863 10553 14897
rect 11629 14863 11641 14897
rect 10541 14851 11641 14863
rect 11987 14801 13087 14813
rect 11987 14767 11999 14801
rect 13075 14767 13087 14801
rect 11987 14755 13087 14767
rect 10541 14639 11641 14651
rect 10541 14605 10553 14639
rect 11629 14605 11641 14639
rect 10541 14593 11641 14605
rect 11987 14583 13087 14595
rect 11987 14549 11999 14583
rect 13075 14549 13087 14583
rect 11987 14537 13087 14549
rect 10541 14473 11641 14485
rect 10541 14439 10553 14473
rect 11629 14439 11641 14473
rect 10541 14427 11641 14439
rect 11987 14441 13087 14453
rect 11987 14407 11999 14441
rect 13075 14407 13087 14441
rect 11987 14395 13087 14407
rect 10541 14215 11641 14227
rect 10541 14181 10553 14215
rect 11629 14181 11641 14215
rect 10541 14169 11641 14181
rect 11987 14223 13087 14235
rect 11987 14189 11999 14223
rect 13075 14189 13087 14223
rect 11987 14177 13087 14189
rect 5930 13855 7030 13867
rect 5930 13821 5942 13855
rect 7018 13821 7030 13855
rect 5930 13809 7030 13821
rect 7406 13811 8506 13823
rect 7406 13777 7418 13811
rect 8494 13777 8506 13811
rect 7406 13765 8506 13777
rect 7406 13673 8506 13685
rect 5930 13637 7030 13649
rect 5930 13603 5942 13637
rect 7018 13603 7030 13637
rect 7406 13639 7418 13673
rect 8494 13639 8506 13673
rect 7406 13627 8506 13639
rect 5930 13591 7030 13603
rect 7406 13513 8506 13525
rect 5930 13495 7030 13507
rect 5930 13461 5942 13495
rect 7018 13461 7030 13495
rect 7406 13479 7418 13513
rect 8494 13479 8506 13513
rect 7406 13467 8506 13479
rect 5930 13449 7030 13461
rect 7406 13375 8506 13387
rect 7406 13341 7418 13375
rect 8494 13341 8506 13375
rect 7406 13329 8506 13341
rect 5930 13277 7030 13289
rect 5930 13243 5942 13277
rect 7018 13243 7030 13277
rect 5930 13231 7030 13243
rect 7376 13231 8476 13243
rect 7376 13197 7388 13231
rect 8464 13197 8476 13231
rect 7376 13185 8476 13197
rect 5930 13135 7030 13147
rect 5930 13101 5942 13135
rect 7018 13101 7030 13135
rect 5930 13089 7030 13101
rect 7376 12973 8476 12985
rect 7376 12939 7388 12973
rect 8464 12939 8476 12973
rect 5930 12917 7030 12929
rect 7376 12927 8476 12939
rect 5930 12883 5942 12917
rect 7018 12883 7030 12917
rect 5930 12871 7030 12883
rect 7376 12807 8476 12819
rect 5930 12775 7030 12787
rect 5930 12741 5942 12775
rect 7018 12741 7030 12775
rect 7376 12773 7388 12807
rect 8464 12773 8476 12807
rect 7376 12761 8476 12773
rect 5930 12729 7030 12741
rect 5930 12557 7030 12569
rect 5930 12523 5942 12557
rect 7018 12523 7030 12557
rect 5930 12511 7030 12523
rect 7376 12549 8476 12561
rect 7376 12515 7388 12549
rect 8464 12515 8476 12549
rect 7376 12503 8476 12515
rect 11987 13855 13087 13867
rect 10511 13811 11611 13823
rect 10511 13777 10523 13811
rect 11599 13777 11611 13811
rect 11987 13821 11999 13855
rect 13075 13821 13087 13855
rect 11987 13809 13087 13821
rect 10511 13765 11611 13777
rect 10511 13673 11611 13685
rect 10511 13639 10523 13673
rect 11599 13639 11611 13673
rect 10511 13627 11611 13639
rect 11987 13637 13087 13649
rect 11987 13603 11999 13637
rect 13075 13603 13087 13637
rect 11987 13591 13087 13603
rect 10511 13513 11611 13525
rect 10511 13479 10523 13513
rect 11599 13479 11611 13513
rect 10511 13467 11611 13479
rect 11987 13495 13087 13507
rect 11987 13461 11999 13495
rect 13075 13461 13087 13495
rect 11987 13449 13087 13461
rect 10511 13375 11611 13387
rect 10511 13341 10523 13375
rect 11599 13341 11611 13375
rect 10511 13329 11611 13341
rect 11987 13277 13087 13289
rect 11987 13243 11999 13277
rect 13075 13243 13087 13277
rect 10541 13231 11641 13243
rect 11987 13231 13087 13243
rect 10541 13197 10553 13231
rect 11629 13197 11641 13231
rect 10541 13185 11641 13197
rect 11987 13135 13087 13147
rect 11987 13101 11999 13135
rect 13075 13101 13087 13135
rect 11987 13089 13087 13101
rect 10541 12973 11641 12985
rect 10541 12939 10553 12973
rect 11629 12939 11641 12973
rect 10541 12927 11641 12939
rect 11987 12917 13087 12929
rect 11987 12883 11999 12917
rect 13075 12883 13087 12917
rect 11987 12871 13087 12883
rect 10541 12807 11641 12819
rect 10541 12773 10553 12807
rect 11629 12773 11641 12807
rect 10541 12761 11641 12773
rect 11987 12775 13087 12787
rect 11987 12741 11999 12775
rect 13075 12741 13087 12775
rect 11987 12729 13087 12741
rect 10541 12549 11641 12561
rect 10541 12515 10553 12549
rect 11629 12515 11641 12549
rect 10541 12503 11641 12515
rect 11987 12557 13087 12569
rect 11987 12523 11999 12557
rect 13075 12523 13087 12557
rect 11987 12511 13087 12523
rect 5930 12189 7030 12201
rect 5930 12155 5942 12189
rect 7018 12155 7030 12189
rect 5930 12143 7030 12155
rect 7406 12145 8506 12157
rect 7406 12111 7418 12145
rect 8494 12111 8506 12145
rect 7406 12099 8506 12111
rect 7406 12007 8506 12019
rect 5930 11971 7030 11983
rect 5930 11937 5942 11971
rect 7018 11937 7030 11971
rect 7406 11973 7418 12007
rect 8494 11973 8506 12007
rect 7406 11961 8506 11973
rect 5930 11925 7030 11937
rect 7406 11847 8506 11859
rect 5930 11829 7030 11841
rect 5930 11795 5942 11829
rect 7018 11795 7030 11829
rect 7406 11813 7418 11847
rect 8494 11813 8506 11847
rect 7406 11801 8506 11813
rect 5930 11783 7030 11795
rect 7406 11709 8506 11721
rect 7406 11675 7418 11709
rect 8494 11675 8506 11709
rect 7406 11663 8506 11675
rect 5930 11611 7030 11623
rect 5930 11577 5942 11611
rect 7018 11577 7030 11611
rect 5930 11565 7030 11577
rect 7376 11565 8476 11577
rect 7376 11531 7388 11565
rect 8464 11531 8476 11565
rect 7376 11519 8476 11531
rect 5930 11469 7030 11481
rect 5930 11435 5942 11469
rect 7018 11435 7030 11469
rect 5930 11423 7030 11435
rect 7376 11307 8476 11319
rect 7376 11273 7388 11307
rect 8464 11273 8476 11307
rect 5930 11251 7030 11263
rect 7376 11261 8476 11273
rect 5930 11217 5942 11251
rect 7018 11217 7030 11251
rect 5930 11205 7030 11217
rect 7376 11141 8476 11153
rect 5930 11109 7030 11121
rect 5930 11075 5942 11109
rect 7018 11075 7030 11109
rect 7376 11107 7388 11141
rect 8464 11107 8476 11141
rect 7376 11095 8476 11107
rect 5930 11063 7030 11075
rect 5930 10891 7030 10903
rect 5930 10857 5942 10891
rect 7018 10857 7030 10891
rect 5930 10845 7030 10857
rect 7376 10883 8476 10895
rect 7376 10849 7388 10883
rect 8464 10849 8476 10883
rect 7376 10837 8476 10849
rect 11987 12189 13087 12201
rect 10511 12145 11611 12157
rect 10511 12111 10523 12145
rect 11599 12111 11611 12145
rect 11987 12155 11999 12189
rect 13075 12155 13087 12189
rect 11987 12143 13087 12155
rect 10511 12099 11611 12111
rect 10511 12007 11611 12019
rect 10511 11973 10523 12007
rect 11599 11973 11611 12007
rect 10511 11961 11611 11973
rect 11987 11971 13087 11983
rect 11987 11937 11999 11971
rect 13075 11937 13087 11971
rect 11987 11925 13087 11937
rect 10511 11847 11611 11859
rect 10511 11813 10523 11847
rect 11599 11813 11611 11847
rect 10511 11801 11611 11813
rect 11987 11829 13087 11841
rect 11987 11795 11999 11829
rect 13075 11795 13087 11829
rect 11987 11783 13087 11795
rect 10511 11709 11611 11721
rect 10511 11675 10523 11709
rect 11599 11675 11611 11709
rect 10511 11663 11611 11675
rect 11987 11611 13087 11623
rect 11987 11577 11999 11611
rect 13075 11577 13087 11611
rect 10541 11565 11641 11577
rect 11987 11565 13087 11577
rect 10541 11531 10553 11565
rect 11629 11531 11641 11565
rect 10541 11519 11641 11531
rect 11987 11469 13087 11481
rect 11987 11435 11999 11469
rect 13075 11435 13087 11469
rect 11987 11423 13087 11435
rect 10541 11307 11641 11319
rect 10541 11273 10553 11307
rect 11629 11273 11641 11307
rect 10541 11261 11641 11273
rect 11987 11251 13087 11263
rect 11987 11217 11999 11251
rect 13075 11217 13087 11251
rect 11987 11205 13087 11217
rect 10541 11141 11641 11153
rect 10541 11107 10553 11141
rect 11629 11107 11641 11141
rect 10541 11095 11641 11107
rect 11987 11109 13087 11121
rect 11987 11075 11999 11109
rect 13075 11075 13087 11109
rect 11987 11063 13087 11075
rect 10541 10883 11641 10895
rect 10541 10849 10553 10883
rect 11629 10849 11641 10883
rect 10541 10837 11641 10849
rect 11987 10891 13087 10903
rect 11987 10857 11999 10891
rect 13075 10857 13087 10891
rect 11987 10845 13087 10857
rect 5930 10523 7030 10535
rect 5930 10489 5942 10523
rect 7018 10489 7030 10523
rect 5930 10477 7030 10489
rect 7406 10479 8506 10491
rect 7406 10445 7418 10479
rect 8494 10445 8506 10479
rect 7406 10433 8506 10445
rect 7406 10341 8506 10353
rect 5930 10305 7030 10317
rect 5930 10271 5942 10305
rect 7018 10271 7030 10305
rect 7406 10307 7418 10341
rect 8494 10307 8506 10341
rect 7406 10295 8506 10307
rect 5930 10259 7030 10271
rect 7406 10181 8506 10193
rect 5930 10163 7030 10175
rect 5930 10129 5942 10163
rect 7018 10129 7030 10163
rect 7406 10147 7418 10181
rect 8494 10147 8506 10181
rect 7406 10135 8506 10147
rect 5930 10117 7030 10129
rect 7406 10043 8506 10055
rect 7406 10009 7418 10043
rect 8494 10009 8506 10043
rect 7406 9997 8506 10009
rect 5930 9945 7030 9957
rect 5930 9911 5942 9945
rect 7018 9911 7030 9945
rect 5930 9899 7030 9911
rect 7376 9899 8476 9911
rect 7376 9865 7388 9899
rect 8464 9865 8476 9899
rect 7376 9853 8476 9865
rect 5930 9803 7030 9815
rect 5930 9769 5942 9803
rect 7018 9769 7030 9803
rect 5930 9757 7030 9769
rect 7376 9641 8476 9653
rect 7376 9607 7388 9641
rect 8464 9607 8476 9641
rect 5930 9585 7030 9597
rect 7376 9595 8476 9607
rect 5930 9551 5942 9585
rect 7018 9551 7030 9585
rect 5930 9539 7030 9551
rect 7376 9475 8476 9487
rect 5930 9443 7030 9455
rect 5930 9409 5942 9443
rect 7018 9409 7030 9443
rect 7376 9441 7388 9475
rect 8464 9441 8476 9475
rect 7376 9429 8476 9441
rect 5930 9397 7030 9409
rect 5930 9225 7030 9237
rect 5930 9191 5942 9225
rect 7018 9191 7030 9225
rect 5930 9179 7030 9191
rect 7376 9217 8476 9229
rect 7376 9183 7388 9217
rect 8464 9183 8476 9217
rect 7376 9171 8476 9183
rect 11987 10523 13087 10535
rect 10511 10479 11611 10491
rect 10511 10445 10523 10479
rect 11599 10445 11611 10479
rect 11987 10489 11999 10523
rect 13075 10489 13087 10523
rect 11987 10477 13087 10489
rect 10511 10433 11611 10445
rect 10511 10341 11611 10353
rect 10511 10307 10523 10341
rect 11599 10307 11611 10341
rect 10511 10295 11611 10307
rect 11987 10305 13087 10317
rect 11987 10271 11999 10305
rect 13075 10271 13087 10305
rect 11987 10259 13087 10271
rect 10511 10181 11611 10193
rect 10511 10147 10523 10181
rect 11599 10147 11611 10181
rect 10511 10135 11611 10147
rect 11987 10163 13087 10175
rect 11987 10129 11999 10163
rect 13075 10129 13087 10163
rect 11987 10117 13087 10129
rect 10511 10043 11611 10055
rect 10511 10009 10523 10043
rect 11599 10009 11611 10043
rect 10511 9997 11611 10009
rect 11987 9945 13087 9957
rect 11987 9911 11999 9945
rect 13075 9911 13087 9945
rect 10541 9899 11641 9911
rect 11987 9899 13087 9911
rect 10541 9865 10553 9899
rect 11629 9865 11641 9899
rect 10541 9853 11641 9865
rect 11987 9803 13087 9815
rect 11987 9769 11999 9803
rect 13075 9769 13087 9803
rect 11987 9757 13087 9769
rect 10541 9641 11641 9653
rect 10541 9607 10553 9641
rect 11629 9607 11641 9641
rect 10541 9595 11641 9607
rect 11987 9585 13087 9597
rect 11987 9551 11999 9585
rect 13075 9551 13087 9585
rect 11987 9539 13087 9551
rect 10541 9475 11641 9487
rect 10541 9441 10553 9475
rect 11629 9441 11641 9475
rect 10541 9429 11641 9441
rect 11987 9443 13087 9455
rect 11987 9409 11999 9443
rect 13075 9409 13087 9443
rect 11987 9397 13087 9409
rect 10541 9217 11641 9229
rect 10541 9183 10553 9217
rect 11629 9183 11641 9217
rect 10541 9171 11641 9183
rect 11987 9225 13087 9237
rect 11987 9191 11999 9225
rect 13075 9191 13087 9225
rect 11987 9179 13087 9191
rect 5930 8857 7030 8869
rect 5930 8823 5942 8857
rect 7018 8823 7030 8857
rect 5930 8811 7030 8823
rect 7406 8813 8506 8825
rect 7406 8779 7418 8813
rect 8494 8779 8506 8813
rect 7406 8767 8506 8779
rect 7406 8675 8506 8687
rect 5930 8639 7030 8651
rect 5930 8605 5942 8639
rect 7018 8605 7030 8639
rect 7406 8641 7418 8675
rect 8494 8641 8506 8675
rect 7406 8629 8506 8641
rect 5930 8593 7030 8605
rect 7406 8515 8506 8527
rect 5930 8497 7030 8509
rect 5930 8463 5942 8497
rect 7018 8463 7030 8497
rect 7406 8481 7418 8515
rect 8494 8481 8506 8515
rect 7406 8469 8506 8481
rect 5930 8451 7030 8463
rect 7406 8377 8506 8389
rect 7406 8343 7418 8377
rect 8494 8343 8506 8377
rect 7406 8331 8506 8343
rect 5930 8279 7030 8291
rect 5930 8245 5942 8279
rect 7018 8245 7030 8279
rect 5930 8233 7030 8245
rect 7376 8233 8476 8245
rect 7376 8199 7388 8233
rect 8464 8199 8476 8233
rect 7376 8187 8476 8199
rect 5930 8137 7030 8149
rect 5930 8103 5942 8137
rect 7018 8103 7030 8137
rect 5930 8091 7030 8103
rect 7376 7975 8476 7987
rect 7376 7941 7388 7975
rect 8464 7941 8476 7975
rect 5930 7919 7030 7931
rect 7376 7929 8476 7941
rect 5930 7885 5942 7919
rect 7018 7885 7030 7919
rect 5930 7873 7030 7885
rect 7376 7809 8476 7821
rect 5930 7777 7030 7789
rect 5930 7743 5942 7777
rect 7018 7743 7030 7777
rect 7376 7775 7388 7809
rect 8464 7775 8476 7809
rect 7376 7763 8476 7775
rect 5930 7731 7030 7743
rect 5930 7559 7030 7571
rect 5930 7525 5942 7559
rect 7018 7525 7030 7559
rect 5930 7513 7030 7525
rect 7376 7551 8476 7563
rect 7376 7517 7388 7551
rect 8464 7517 8476 7551
rect 7376 7505 8476 7517
rect 11987 8857 13087 8869
rect 10511 8813 11611 8825
rect 10511 8779 10523 8813
rect 11599 8779 11611 8813
rect 11987 8823 11999 8857
rect 13075 8823 13087 8857
rect 11987 8811 13087 8823
rect 10511 8767 11611 8779
rect 10511 8675 11611 8687
rect 10511 8641 10523 8675
rect 11599 8641 11611 8675
rect 10511 8629 11611 8641
rect 11987 8639 13087 8651
rect 11987 8605 11999 8639
rect 13075 8605 13087 8639
rect 11987 8593 13087 8605
rect 10511 8515 11611 8527
rect 10511 8481 10523 8515
rect 11599 8481 11611 8515
rect 10511 8469 11611 8481
rect 11987 8497 13087 8509
rect 11987 8463 11999 8497
rect 13075 8463 13087 8497
rect 11987 8451 13087 8463
rect 10511 8377 11611 8389
rect 10511 8343 10523 8377
rect 11599 8343 11611 8377
rect 10511 8331 11611 8343
rect 11987 8279 13087 8291
rect 11987 8245 11999 8279
rect 13075 8245 13087 8279
rect 10541 8233 11641 8245
rect 11987 8233 13087 8245
rect 10541 8199 10553 8233
rect 11629 8199 11641 8233
rect 10541 8187 11641 8199
rect 11987 8137 13087 8149
rect 11987 8103 11999 8137
rect 13075 8103 13087 8137
rect 11987 8091 13087 8103
rect 10541 7975 11641 7987
rect 10541 7941 10553 7975
rect 11629 7941 11641 7975
rect 10541 7929 11641 7941
rect 11987 7919 13087 7931
rect 11987 7885 11999 7919
rect 13075 7885 13087 7919
rect 11987 7873 13087 7885
rect 10541 7809 11641 7821
rect 10541 7775 10553 7809
rect 11629 7775 11641 7809
rect 10541 7763 11641 7775
rect 11987 7777 13087 7789
rect 11987 7743 11999 7777
rect 13075 7743 13087 7777
rect 11987 7731 13087 7743
rect 10541 7551 11641 7563
rect 10541 7517 10553 7551
rect 11629 7517 11641 7551
rect 10541 7505 11641 7517
rect 11987 7559 13087 7571
rect 11987 7525 11999 7559
rect 13075 7525 13087 7559
rect 11987 7513 13087 7525
rect 16238 17496 17438 17508
rect 16238 17462 16250 17496
rect 17426 17462 17438 17496
rect 16238 17450 17438 17462
rect 16238 17260 17438 17272
rect 16238 17226 16250 17260
rect 17426 17226 17438 17260
rect 16238 17214 17438 17226
rect 16238 17126 17438 17138
rect 16238 17092 16250 17126
rect 17426 17092 17438 17126
rect 16238 17080 17438 17092
rect 16238 16890 17438 16902
rect 16238 16856 16250 16890
rect 17426 16856 17438 16890
rect 16238 16844 17438 16856
rect 16474 16644 16532 16656
rect 16474 16324 16486 16644
rect 16520 16324 16532 16644
rect 16474 16312 16532 16324
rect 17152 16644 17210 16656
rect 17152 16324 17164 16644
rect 17198 16324 17210 16644
rect 17362 16572 17420 16584
rect 17362 16432 17374 16572
rect 17408 16432 17420 16572
rect 17362 16420 17420 16432
rect 17630 16572 17688 16584
rect 17630 16432 17642 16572
rect 17676 16432 17688 16572
rect 17630 16420 17688 16432
rect 17152 16312 17210 16324
rect 14490 11662 14548 11674
rect 14490 10648 14502 11662
rect 14536 10648 14548 11662
rect 14490 10636 14548 10648
rect 14834 11662 14892 11674
rect 14834 10648 14846 11662
rect 14880 10648 14892 11662
rect 14834 10636 14892 10648
rect 14490 10406 14548 10418
rect 14490 9392 14502 10406
rect 14536 9392 14548 10406
rect 14490 9380 14548 9392
rect 14834 10406 14892 10418
rect 14834 9392 14846 10406
rect 14880 9392 14892 10406
rect 14834 9380 14892 9392
rect 14464 8586 14522 8598
rect 14464 7590 14476 8586
rect 14510 7590 14522 8586
rect 14464 7578 14522 7590
rect 14654 8586 14712 8598
rect 14654 7590 14666 8586
rect 14700 7590 14712 8586
rect 14654 7578 14712 7590
rect 14864 8586 14922 8598
rect 14864 7590 14876 8586
rect 14910 7590 14922 8586
rect 14864 7578 14922 7590
rect 15054 8586 15112 8598
rect 15054 7590 15066 8586
rect 15100 7590 15112 8586
rect 15054 7578 15112 7590
rect 15264 8586 15322 8598
rect 15264 7590 15276 8586
rect 15310 7590 15322 8586
rect 15264 7578 15322 7590
rect 15454 8586 15512 8598
rect 15454 7590 15466 8586
rect 15500 7590 15512 8586
rect 15454 7578 15512 7590
rect 15664 8586 15722 8598
rect 15664 7590 15676 8586
rect 15710 7590 15722 8586
rect 15664 7578 15722 7590
rect 15854 8586 15912 8598
rect 15854 7590 15866 8586
rect 15900 7590 15912 8586
rect 15854 7578 15912 7590
rect 16064 8586 16122 8598
rect 16064 7590 16076 8586
rect 16110 7590 16122 8586
rect 16064 7578 16122 7590
rect 16254 8586 16312 8598
rect 16254 7590 16266 8586
rect 16300 7590 16312 8586
rect 16254 7578 16312 7590
rect 16464 8586 16522 8598
rect 16464 7590 16476 8586
rect 16510 7590 16522 8586
rect 16464 7578 16522 7590
rect 16654 8586 16712 8598
rect 16654 7590 16666 8586
rect 16700 7590 16712 8586
rect 16654 7578 16712 7590
rect 16864 8586 16922 8598
rect 16864 7590 16876 8586
rect 16910 7590 16922 8586
rect 16864 7578 16922 7590
rect 17054 8586 17112 8598
rect 17054 7590 17066 8586
rect 17100 7590 17112 8586
rect 17054 7578 17112 7590
rect 17264 8586 17322 8598
rect 17264 7590 17276 8586
rect 17310 7590 17322 8586
rect 17264 7578 17322 7590
rect 17454 8586 17512 8598
rect 17454 7590 17466 8586
rect 17500 7590 17512 8586
rect 17454 7578 17512 7590
rect 17664 8586 17722 8598
rect 17664 7590 17676 8586
rect 17710 7590 17722 8586
rect 17664 7578 17722 7590
rect 17854 8586 17912 8598
rect 17854 7590 17866 8586
rect 17900 7590 17912 8586
rect 17854 7578 17912 7590
rect 18064 8586 18122 8598
rect 18064 7590 18076 8586
rect 18110 7590 18122 8586
rect 18064 7578 18122 7590
rect 18254 8586 18312 8598
rect 18254 7590 18266 8586
rect 18300 7590 18312 8586
rect 18254 7578 18312 7590
<< pdiff >>
rect 1328 19186 1386 19198
rect 1328 19110 1340 19186
rect 1374 19110 1386 19186
rect 1328 19098 1386 19110
rect 1786 19186 1844 19198
rect 1786 19110 1798 19186
rect 1832 19110 1844 19186
rect 1786 19098 1844 19110
rect 2028 19186 2086 19198
rect 2028 19110 2040 19186
rect 2074 19110 2086 19186
rect 2028 19098 2086 19110
rect 2486 19186 2544 19198
rect 2486 19110 2498 19186
rect 2532 19110 2544 19186
rect 2486 19098 2544 19110
rect 1328 18802 1386 18814
rect 1328 18326 1340 18802
rect 1374 18326 1386 18802
rect 1328 18314 1386 18326
rect 1786 18802 1844 18814
rect 1786 18326 1798 18802
rect 1832 18326 1844 18802
rect 1786 18314 1844 18326
rect 2028 18802 2086 18814
rect 2028 18326 2040 18802
rect 2074 18326 2086 18802
rect 2028 18314 2086 18326
rect 2486 18802 2544 18814
rect 2486 18326 2498 18802
rect 2532 18326 2544 18802
rect 2486 18314 2544 18326
rect 1328 18018 1386 18030
rect 1328 17542 1340 18018
rect 1374 17542 1386 18018
rect 1328 17530 1386 17542
rect 1786 18018 1844 18030
rect 1786 17542 1798 18018
rect 1832 17542 1844 18018
rect 1786 17530 1844 17542
rect 2028 18018 2086 18030
rect 2028 17542 2040 18018
rect 2074 17542 2086 18018
rect 2028 17530 2086 17542
rect 2486 18018 2544 18030
rect 2486 17542 2498 18018
rect 2532 17542 2544 18018
rect 2486 17530 2544 17542
rect 1328 17234 1386 17246
rect 1328 16758 1340 17234
rect 1374 16758 1386 17234
rect 1328 16746 1386 16758
rect 1786 17234 1844 17246
rect 1786 16758 1798 17234
rect 1832 16758 1844 17234
rect 1786 16746 1844 16758
rect 2028 17234 2086 17246
rect 2028 16758 2040 17234
rect 2074 16758 2086 17234
rect 2028 16746 2086 16758
rect 2486 17234 2544 17246
rect 2486 16758 2498 17234
rect 2532 16758 2544 17234
rect 2486 16746 2544 16758
rect 1328 16450 1386 16462
rect 1328 15974 1340 16450
rect 1374 15974 1386 16450
rect 1328 15962 1386 15974
rect 1786 16450 1844 16462
rect 1786 15974 1798 16450
rect 1832 15974 1844 16450
rect 1786 15962 1844 15974
rect 2028 16450 2086 16462
rect 2028 15974 2040 16450
rect 2074 15974 2086 16450
rect 2028 15962 2086 15974
rect 2486 16450 2544 16462
rect 2486 15974 2498 16450
rect 2532 15974 2544 16450
rect 2486 15962 2544 15974
rect 1328 15666 1386 15678
rect 1328 15590 1340 15666
rect 1374 15590 1386 15666
rect 1328 15578 1386 15590
rect 1786 15666 1844 15678
rect 1786 15590 1798 15666
rect 1832 15590 1844 15666
rect 1786 15578 1844 15590
rect 2028 15666 2086 15678
rect 2028 15590 2040 15666
rect 2074 15590 2086 15666
rect 2028 15578 2086 15590
rect 2486 15666 2544 15678
rect 2486 15590 2498 15666
rect 2532 15590 2544 15666
rect 2486 15578 2544 15590
rect -163 12726 237 12738
rect -163 12692 -151 12726
rect 225 12692 237 12726
rect -163 12680 237 12692
rect 473 12726 873 12738
rect 473 12692 485 12726
rect 861 12692 873 12726
rect 473 12680 873 12692
rect 1109 12726 1509 12738
rect 1109 12692 1121 12726
rect 1497 12692 1509 12726
rect 1109 12680 1509 12692
rect 1745 12726 2145 12738
rect 1745 12692 1757 12726
rect 2133 12692 2145 12726
rect 1745 12680 2145 12692
rect -163 12568 237 12580
rect -163 12534 -151 12568
rect 225 12534 237 12568
rect -163 12522 237 12534
rect 473 12568 873 12580
rect 473 12534 485 12568
rect 861 12534 873 12568
rect 473 12522 873 12534
rect 1109 12568 1509 12580
rect 1109 12534 1121 12568
rect 1497 12534 1509 12568
rect 1109 12522 1509 12534
rect 1745 12568 2145 12580
rect 1745 12534 1757 12568
rect 2133 12534 2145 12568
rect 1745 12522 2145 12534
rect 721 11887 779 11899
rect 721 11735 733 11887
rect 767 11735 779 11887
rect 721 11723 779 11735
rect 2173 11887 2231 11899
rect 2173 11735 2185 11887
rect 2219 11735 2231 11887
rect 2173 11723 2231 11735
rect 343 10985 401 10997
rect 343 10323 355 10985
rect 389 10323 401 10985
rect 343 10311 401 10323
rect 955 10985 1013 10997
rect 955 10323 967 10985
rect 1001 10323 1013 10985
rect 1337 10979 1395 10991
rect 1337 10903 1349 10979
rect 1383 10903 1395 10979
rect 1337 10891 1395 10903
rect 2195 10979 2253 10991
rect 2195 10903 2207 10979
rect 2241 10903 2253 10979
rect 2195 10891 2253 10903
rect 955 10311 1013 10323
rect 1263 10587 1321 10599
rect 1263 10137 1275 10587
rect 1309 10137 1321 10587
rect 1263 10125 1321 10137
rect 2197 10587 2255 10599
rect 2197 10137 2209 10587
rect 2243 10137 2255 10587
rect 2197 10125 2255 10137
rect 1097 9240 1155 9252
rect 1097 8764 1109 9240
rect 1143 8764 1155 9240
rect 1097 8752 1155 8764
rect 1555 9240 1613 9252
rect 1555 8764 1567 9240
rect 1601 8764 1613 9240
rect 1555 8752 1613 8764
rect 1797 9240 1855 9252
rect 1797 8764 1809 9240
rect 1843 8764 1855 9240
rect 1797 8752 1855 8764
rect 2255 9240 2313 9252
rect 2255 8764 2267 9240
rect 2301 8764 2313 9240
rect 2255 8752 2313 8764
rect 1097 8456 1155 8468
rect 1097 7980 1109 8456
rect 1143 7980 1155 8456
rect 1097 7968 1155 7980
rect 1555 8456 1613 8468
rect 1555 7980 1567 8456
rect 1601 7980 1613 8456
rect 1555 7968 1613 7980
rect 1797 8456 1855 8468
rect 1797 7980 1809 8456
rect 1843 7980 1855 8456
rect 1797 7968 1855 7980
rect 2255 8456 2313 8468
rect 2255 7980 2267 8456
rect 2301 7980 2313 8456
rect 2255 7968 2313 7980
rect 3024 19202 3082 19214
rect 3024 19126 3036 19202
rect 3070 19126 3082 19202
rect 3024 19114 3082 19126
rect 3482 19202 3540 19214
rect 3482 19126 3494 19202
rect 3528 19126 3540 19202
rect 3482 19114 3540 19126
rect 3724 19202 3782 19214
rect 3724 19126 3736 19202
rect 3770 19126 3782 19202
rect 3724 19114 3782 19126
rect 4182 19202 4240 19214
rect 4182 19126 4194 19202
rect 4228 19126 4240 19202
rect 4182 19114 4240 19126
rect 3024 18818 3082 18830
rect 3024 18342 3036 18818
rect 3070 18342 3082 18818
rect 3024 18330 3082 18342
rect 3482 18818 3540 18830
rect 3482 18342 3494 18818
rect 3528 18342 3540 18818
rect 3482 18330 3540 18342
rect 3724 18818 3782 18830
rect 3724 18342 3736 18818
rect 3770 18342 3782 18818
rect 3724 18330 3782 18342
rect 4182 18818 4240 18830
rect 4182 18342 4194 18818
rect 4228 18342 4240 18818
rect 4182 18330 4240 18342
rect 3024 18034 3082 18046
rect 3024 17558 3036 18034
rect 3070 17558 3082 18034
rect 3024 17546 3082 17558
rect 3482 18034 3540 18046
rect 3482 17558 3494 18034
rect 3528 17558 3540 18034
rect 3482 17546 3540 17558
rect 3724 18034 3782 18046
rect 3724 17558 3736 18034
rect 3770 17558 3782 18034
rect 3724 17546 3782 17558
rect 4182 18034 4240 18046
rect 4182 17558 4194 18034
rect 4228 17558 4240 18034
rect 4182 17546 4240 17558
rect 3024 17250 3082 17262
rect 3024 16774 3036 17250
rect 3070 16774 3082 17250
rect 3024 16762 3082 16774
rect 3482 17250 3540 17262
rect 3482 16774 3494 17250
rect 3528 16774 3540 17250
rect 3482 16762 3540 16774
rect 3724 17250 3782 17262
rect 3724 16774 3736 17250
rect 3770 16774 3782 17250
rect 3724 16762 3782 16774
rect 4182 17250 4240 17262
rect 4182 16774 4194 17250
rect 4228 16774 4240 17250
rect 4182 16762 4240 16774
rect 3024 16466 3082 16478
rect 3024 15990 3036 16466
rect 3070 15990 3082 16466
rect 3024 15978 3082 15990
rect 3482 16466 3540 16478
rect 3482 15990 3494 16466
rect 3528 15990 3540 16466
rect 3482 15978 3540 15990
rect 3724 16466 3782 16478
rect 3724 15990 3736 16466
rect 3770 15990 3782 16466
rect 3724 15978 3782 15990
rect 4182 16466 4240 16478
rect 4182 15990 4194 16466
rect 4228 15990 4240 16466
rect 4182 15978 4240 15990
rect 3024 15682 3082 15694
rect 3024 15206 3036 15682
rect 3070 15206 3082 15682
rect 3024 15194 3082 15206
rect 3482 15682 3540 15694
rect 3482 15206 3494 15682
rect 3528 15206 3540 15682
rect 3482 15194 3540 15206
rect 3724 15682 3782 15694
rect 3724 15206 3736 15682
rect 3770 15206 3782 15682
rect 3724 15194 3782 15206
rect 4182 15682 4240 15694
rect 4182 15206 4194 15682
rect 4228 15206 4240 15682
rect 4182 15194 4240 15206
rect 3024 14898 3082 14910
rect 3024 14422 3036 14898
rect 3070 14422 3082 14898
rect 3024 14410 3082 14422
rect 3482 14898 3540 14910
rect 3482 14422 3494 14898
rect 3528 14422 3540 14898
rect 3482 14410 3540 14422
rect 3724 14898 3782 14910
rect 3724 14422 3736 14898
rect 3770 14422 3782 14898
rect 3724 14410 3782 14422
rect 4182 14898 4240 14910
rect 4182 14422 4194 14898
rect 4228 14422 4240 14898
rect 4182 14410 4240 14422
rect 3024 14114 3082 14126
rect 3024 13638 3036 14114
rect 3070 13638 3082 14114
rect 3024 13626 3082 13638
rect 3482 14114 3540 14126
rect 3482 13638 3494 14114
rect 3528 13638 3540 14114
rect 3482 13626 3540 13638
rect 3724 14114 3782 14126
rect 3724 13638 3736 14114
rect 3770 13638 3782 14114
rect 3724 13626 3782 13638
rect 4182 14114 4240 14126
rect 4182 13638 4194 14114
rect 4228 13638 4240 14114
rect 4182 13626 4240 13638
rect 3024 13330 3082 13342
rect 3024 12854 3036 13330
rect 3070 12854 3082 13330
rect 3024 12842 3082 12854
rect 3482 13330 3540 13342
rect 3482 12854 3494 13330
rect 3528 12854 3540 13330
rect 3482 12842 3540 12854
rect 3724 13330 3782 13342
rect 3724 12854 3736 13330
rect 3770 12854 3782 13330
rect 3724 12842 3782 12854
rect 4182 13330 4240 13342
rect 4182 12854 4194 13330
rect 4228 12854 4240 13330
rect 4182 12842 4240 12854
rect 3024 12546 3082 12558
rect 3024 12070 3036 12546
rect 3070 12070 3082 12546
rect 3024 12058 3082 12070
rect 3482 12546 3540 12558
rect 3482 12070 3494 12546
rect 3528 12070 3540 12546
rect 3482 12058 3540 12070
rect 3724 12546 3782 12558
rect 3724 12070 3736 12546
rect 3770 12070 3782 12546
rect 3724 12058 3782 12070
rect 4182 12546 4240 12558
rect 4182 12070 4194 12546
rect 4228 12070 4240 12546
rect 4182 12058 4240 12070
rect 3024 11762 3082 11774
rect 3024 11286 3036 11762
rect 3070 11286 3082 11762
rect 3024 11274 3082 11286
rect 3482 11762 3540 11774
rect 3482 11286 3494 11762
rect 3528 11286 3540 11762
rect 3482 11274 3540 11286
rect 3724 11762 3782 11774
rect 3724 11286 3736 11762
rect 3770 11286 3782 11762
rect 3724 11274 3782 11286
rect 4182 11762 4240 11774
rect 4182 11286 4194 11762
rect 4228 11286 4240 11762
rect 4182 11274 4240 11286
rect 3024 10978 3082 10990
rect 3024 10502 3036 10978
rect 3070 10502 3082 10978
rect 3024 10490 3082 10502
rect 3482 10978 3540 10990
rect 3482 10502 3494 10978
rect 3528 10502 3540 10978
rect 3482 10490 3540 10502
rect 3724 10978 3782 10990
rect 3724 10502 3736 10978
rect 3770 10502 3782 10978
rect 3724 10490 3782 10502
rect 4182 10978 4240 10990
rect 4182 10502 4194 10978
rect 4228 10502 4240 10978
rect 4182 10490 4240 10502
rect 3024 10194 3082 10206
rect 3024 9718 3036 10194
rect 3070 9718 3082 10194
rect 3024 9706 3082 9718
rect 3482 10194 3540 10206
rect 3482 9718 3494 10194
rect 3528 9718 3540 10194
rect 3482 9706 3540 9718
rect 3724 10194 3782 10206
rect 3724 9718 3736 10194
rect 3770 9718 3782 10194
rect 3724 9706 3782 9718
rect 4182 10194 4240 10206
rect 4182 9718 4194 10194
rect 4228 9718 4240 10194
rect 4182 9706 4240 9718
rect 3024 9410 3082 9422
rect 3024 8934 3036 9410
rect 3070 8934 3082 9410
rect 3024 8922 3082 8934
rect 3482 9410 3540 9422
rect 3482 8934 3494 9410
rect 3528 8934 3540 9410
rect 3482 8922 3540 8934
rect 3724 9410 3782 9422
rect 3724 8934 3736 9410
rect 3770 8934 3782 9410
rect 3724 8922 3782 8934
rect 4182 9410 4240 9422
rect 4182 8934 4194 9410
rect 4228 8934 4240 9410
rect 4182 8922 4240 8934
rect 3024 8626 3082 8638
rect 3024 8150 3036 8626
rect 3070 8150 3082 8626
rect 3024 8138 3082 8150
rect 3482 8626 3540 8638
rect 3482 8150 3494 8626
rect 3528 8150 3540 8626
rect 3482 8138 3540 8150
rect 3724 8626 3782 8638
rect 3724 8150 3736 8626
rect 3770 8150 3782 8626
rect 3724 8138 3782 8150
rect 4182 8626 4240 8638
rect 4182 8150 4194 8626
rect 4228 8150 4240 8626
rect 4182 8138 4240 8150
rect 3024 7842 3082 7854
rect 3024 7766 3036 7842
rect 3070 7766 3082 7842
rect 3024 7754 3082 7766
rect 3482 7842 3540 7854
rect 3482 7766 3494 7842
rect 3528 7766 3540 7842
rect 3482 7754 3540 7766
rect 3724 7842 3782 7854
rect 3724 7766 3736 7842
rect 3770 7766 3782 7842
rect 3724 7754 3782 7766
rect 4182 7842 4240 7854
rect 4182 7766 4194 7842
rect 4228 7766 4240 7842
rect 4182 7754 4240 7766
rect 9356 17302 9414 17314
rect 9356 17126 9368 17302
rect 9402 17126 9414 17302
rect 9356 17114 9414 17126
rect 9574 17302 9632 17314
rect 9574 17126 9586 17302
rect 9620 17126 9632 17302
rect 9574 17114 9632 17126
rect 9756 17302 9814 17314
rect 9756 17126 9768 17302
rect 9802 17126 9814 17302
rect 9756 17114 9814 17126
rect 9974 17302 10032 17314
rect 9974 17126 9986 17302
rect 10020 17126 10032 17302
rect 9974 17114 10032 17126
rect 10615 17273 10673 17285
rect 10615 17097 10627 17273
rect 10661 17097 10673 17273
rect 10615 17085 10673 17097
rect 10833 17273 10891 17285
rect 10833 17097 10845 17273
rect 10879 17097 10891 17273
rect 10833 17085 10891 17097
rect 11015 17273 11073 17285
rect 11015 17097 11027 17273
rect 11061 17097 11073 17273
rect 11015 17085 11073 17097
rect 11233 17273 11291 17285
rect 11233 17097 11245 17273
rect 11279 17097 11291 17273
rect 11233 17085 11291 17097
rect 11415 17273 11473 17285
rect 11415 17097 11427 17273
rect 11461 17097 11473 17273
rect 11415 17085 11473 17097
rect 11633 17273 11691 17285
rect 11633 17097 11645 17273
rect 11679 17097 11691 17273
rect 11633 17085 11691 17097
rect 11815 17273 11873 17285
rect 11815 17097 11827 17273
rect 11861 17097 11873 17273
rect 11815 17085 11873 17097
rect 12033 17273 12091 17285
rect 12033 17097 12045 17273
rect 12079 17097 12091 17273
rect 12033 17085 12091 17097
rect 9063 15552 9263 15564
rect 9063 15518 9075 15552
rect 9251 15518 9263 15552
rect 9063 15506 9263 15518
rect 9063 15334 9263 15346
rect 9063 15300 9075 15334
rect 9251 15300 9263 15334
rect 9063 15288 9263 15300
rect 9063 15144 9263 15156
rect 9063 15110 9075 15144
rect 9251 15110 9263 15144
rect 9063 15098 9263 15110
rect 9063 14926 9263 14938
rect 9063 14892 9075 14926
rect 9251 14892 9263 14926
rect 9063 14880 9263 14892
rect 9063 14698 9263 14710
rect 9063 14664 9075 14698
rect 9251 14664 9263 14698
rect 9063 14652 9263 14664
rect 9063 14240 9263 14252
rect 9063 14206 9075 14240
rect 9251 14206 9263 14240
rect 9063 14194 9263 14206
rect 9754 15552 9954 15564
rect 9754 15518 9766 15552
rect 9942 15518 9954 15552
rect 9754 15506 9954 15518
rect 9754 15334 9954 15346
rect 9754 15300 9766 15334
rect 9942 15300 9954 15334
rect 9754 15288 9954 15300
rect 9754 15144 9954 15156
rect 9754 15110 9766 15144
rect 9942 15110 9954 15144
rect 9754 15098 9954 15110
rect 9754 14926 9954 14938
rect 9754 14892 9766 14926
rect 9942 14892 9954 14926
rect 9754 14880 9954 14892
rect 9754 14698 9954 14710
rect 9754 14664 9766 14698
rect 9942 14664 9954 14698
rect 9754 14652 9954 14664
rect 9754 14240 9954 14252
rect 9754 14206 9766 14240
rect 9942 14206 9954 14240
rect 9754 14194 9954 14206
rect 9063 13886 9263 13898
rect 9063 13852 9075 13886
rect 9251 13852 9263 13886
rect 9063 13840 9263 13852
rect 9063 13668 9263 13680
rect 9063 13634 9075 13668
rect 9251 13634 9263 13668
rect 9063 13622 9263 13634
rect 9063 13478 9263 13490
rect 9063 13444 9075 13478
rect 9251 13444 9263 13478
rect 9063 13432 9263 13444
rect 9063 13260 9263 13272
rect 9063 13226 9075 13260
rect 9251 13226 9263 13260
rect 9063 13214 9263 13226
rect 9063 13032 9263 13044
rect 9063 12998 9075 13032
rect 9251 12998 9263 13032
rect 9063 12986 9263 12998
rect 9063 12574 9263 12586
rect 9063 12540 9075 12574
rect 9251 12540 9263 12574
rect 9063 12528 9263 12540
rect 9754 13886 9954 13898
rect 9754 13852 9766 13886
rect 9942 13852 9954 13886
rect 9754 13840 9954 13852
rect 9754 13668 9954 13680
rect 9754 13634 9766 13668
rect 9942 13634 9954 13668
rect 9754 13622 9954 13634
rect 9754 13478 9954 13490
rect 9754 13444 9766 13478
rect 9942 13444 9954 13478
rect 9754 13432 9954 13444
rect 9754 13260 9954 13272
rect 9754 13226 9766 13260
rect 9942 13226 9954 13260
rect 9754 13214 9954 13226
rect 9754 13032 9954 13044
rect 9754 12998 9766 13032
rect 9942 12998 9954 13032
rect 9754 12986 9954 12998
rect 9754 12574 9954 12586
rect 9754 12540 9766 12574
rect 9942 12540 9954 12574
rect 9754 12528 9954 12540
rect 9063 12220 9263 12232
rect 9063 12186 9075 12220
rect 9251 12186 9263 12220
rect 9063 12174 9263 12186
rect 9063 12002 9263 12014
rect 9063 11968 9075 12002
rect 9251 11968 9263 12002
rect 9063 11956 9263 11968
rect 9063 11812 9263 11824
rect 9063 11778 9075 11812
rect 9251 11778 9263 11812
rect 9063 11766 9263 11778
rect 9063 11594 9263 11606
rect 9063 11560 9075 11594
rect 9251 11560 9263 11594
rect 9063 11548 9263 11560
rect 9063 11366 9263 11378
rect 9063 11332 9075 11366
rect 9251 11332 9263 11366
rect 9063 11320 9263 11332
rect 9063 10908 9263 10920
rect 9063 10874 9075 10908
rect 9251 10874 9263 10908
rect 9063 10862 9263 10874
rect 9754 12220 9954 12232
rect 9754 12186 9766 12220
rect 9942 12186 9954 12220
rect 9754 12174 9954 12186
rect 9754 12002 9954 12014
rect 9754 11968 9766 12002
rect 9942 11968 9954 12002
rect 9754 11956 9954 11968
rect 9754 11812 9954 11824
rect 9754 11778 9766 11812
rect 9942 11778 9954 11812
rect 9754 11766 9954 11778
rect 9754 11594 9954 11606
rect 9754 11560 9766 11594
rect 9942 11560 9954 11594
rect 9754 11548 9954 11560
rect 9754 11366 9954 11378
rect 9754 11332 9766 11366
rect 9942 11332 9954 11366
rect 9754 11320 9954 11332
rect 9754 10908 9954 10920
rect 9754 10874 9766 10908
rect 9942 10874 9954 10908
rect 9754 10862 9954 10874
rect 9063 10554 9263 10566
rect 9063 10520 9075 10554
rect 9251 10520 9263 10554
rect 9063 10508 9263 10520
rect 9063 10336 9263 10348
rect 9063 10302 9075 10336
rect 9251 10302 9263 10336
rect 9063 10290 9263 10302
rect 9063 10146 9263 10158
rect 9063 10112 9075 10146
rect 9251 10112 9263 10146
rect 9063 10100 9263 10112
rect 9063 9928 9263 9940
rect 9063 9894 9075 9928
rect 9251 9894 9263 9928
rect 9063 9882 9263 9894
rect 9063 9700 9263 9712
rect 9063 9666 9075 9700
rect 9251 9666 9263 9700
rect 9063 9654 9263 9666
rect 9063 9242 9263 9254
rect 9063 9208 9075 9242
rect 9251 9208 9263 9242
rect 9063 9196 9263 9208
rect 9754 10554 9954 10566
rect 9754 10520 9766 10554
rect 9942 10520 9954 10554
rect 9754 10508 9954 10520
rect 9754 10336 9954 10348
rect 9754 10302 9766 10336
rect 9942 10302 9954 10336
rect 9754 10290 9954 10302
rect 9754 10146 9954 10158
rect 9754 10112 9766 10146
rect 9942 10112 9954 10146
rect 9754 10100 9954 10112
rect 9754 9928 9954 9940
rect 9754 9894 9766 9928
rect 9942 9894 9954 9928
rect 9754 9882 9954 9894
rect 9754 9700 9954 9712
rect 9754 9666 9766 9700
rect 9942 9666 9954 9700
rect 9754 9654 9954 9666
rect 9754 9242 9954 9254
rect 9754 9208 9766 9242
rect 9942 9208 9954 9242
rect 9754 9196 9954 9208
rect 9063 8888 9263 8900
rect 9063 8854 9075 8888
rect 9251 8854 9263 8888
rect 9063 8842 9263 8854
rect 9063 8670 9263 8682
rect 9063 8636 9075 8670
rect 9251 8636 9263 8670
rect 9063 8624 9263 8636
rect 9063 8480 9263 8492
rect 9063 8446 9075 8480
rect 9251 8446 9263 8480
rect 9063 8434 9263 8446
rect 9063 8262 9263 8274
rect 9063 8228 9075 8262
rect 9251 8228 9263 8262
rect 9063 8216 9263 8228
rect 9063 8034 9263 8046
rect 9063 8000 9075 8034
rect 9251 8000 9263 8034
rect 9063 7988 9263 8000
rect 9063 7576 9263 7588
rect 9063 7542 9075 7576
rect 9251 7542 9263 7576
rect 9063 7530 9263 7542
rect 9754 8888 9954 8900
rect 9754 8854 9766 8888
rect 9942 8854 9954 8888
rect 9754 8842 9954 8854
rect 9754 8670 9954 8682
rect 9754 8636 9766 8670
rect 9942 8636 9954 8670
rect 9754 8624 9954 8636
rect 9754 8480 9954 8492
rect 9754 8446 9766 8480
rect 9942 8446 9954 8480
rect 9754 8434 9954 8446
rect 9754 8262 9954 8274
rect 9754 8228 9766 8262
rect 9942 8228 9954 8262
rect 9754 8216 9954 8228
rect 9754 8034 9954 8046
rect 9754 8000 9766 8034
rect 9942 8000 9954 8034
rect 9754 7988 9954 8000
rect 9754 7576 9954 7588
rect 9754 7542 9766 7576
rect 9942 7542 9954 7576
rect 9754 7530 9954 7542
rect 14901 17673 15101 17685
rect 14901 15977 15055 17673
rect 15089 15977 15101 17673
rect 14901 15965 15101 15977
rect 15171 17673 15371 17685
rect 15171 15977 15183 17673
rect 15217 15977 15371 17673
rect 15171 15965 15371 15977
rect 14982 13502 15160 13514
rect 14982 13468 14994 13502
rect 15148 13468 15160 13502
rect 14982 13456 15160 13468
rect 15482 13502 15660 13514
rect 15482 13468 15494 13502
rect 15648 13468 15660 13502
rect 15482 13456 15660 13468
rect 15982 13502 16160 13514
rect 15982 13468 15994 13502
rect 16148 13468 16160 13502
rect 15982 13456 16160 13468
rect 16482 13502 16660 13514
rect 16482 13468 16494 13502
rect 16648 13468 16660 13502
rect 16482 13456 16660 13468
rect 16982 13502 17160 13514
rect 16982 13468 16994 13502
rect 17148 13468 17160 13502
rect 16982 13456 17160 13468
rect 17482 13502 17660 13514
rect 17482 13468 17494 13502
rect 17648 13468 17660 13502
rect 17482 13456 17660 13468
rect 14982 12666 15160 12678
rect 14982 12632 14994 12666
rect 15148 12632 15160 12666
rect 14982 12620 15160 12632
rect 15482 12666 15660 12678
rect 15482 12632 15494 12666
rect 15648 12632 15660 12666
rect 15482 12620 15660 12632
rect 15982 12666 16160 12678
rect 15982 12632 15994 12666
rect 16148 12632 16160 12666
rect 15982 12620 16160 12632
rect 16482 12666 16660 12678
rect 16482 12632 16494 12666
rect 16648 12632 16660 12666
rect 16482 12620 16660 12632
rect 16982 12666 17160 12678
rect 16982 12632 16994 12666
rect 17148 12632 17160 12666
rect 16982 12620 17160 12632
rect 17482 12666 17660 12678
rect 17482 12632 17494 12666
rect 17648 12632 17660 12666
rect 17482 12620 17660 12632
rect 17086 11347 18120 11359
rect 17086 11313 17098 11347
rect 18108 11313 18120 11347
rect 17086 11301 18120 11313
rect 17086 11215 18120 11227
rect 17086 11181 17098 11215
rect 18108 11181 18120 11215
rect 17086 11169 18120 11181
rect 17029 10280 18243 10292
rect 17029 10246 17041 10280
rect 18231 10246 18243 10280
rect 17029 10234 18243 10246
rect 17029 9968 18243 9980
rect 17029 9934 17041 9968
rect 18231 9934 18243 9968
rect 17029 9922 18243 9934
rect 17029 9680 18243 9692
rect 17029 9646 17041 9680
rect 18231 9646 18243 9680
rect 17029 9634 18243 9646
rect 17029 9368 18243 9380
rect 17029 9334 17041 9368
rect 18231 9334 18243 9368
rect 17029 9322 18243 9334
<< ndiffc >>
rect -69 18995 407 19029
rect -69 18737 407 18771
rect -69 18579 407 18613
rect -69 18321 407 18355
rect -69 18163 407 18197
rect -69 17905 407 17939
rect -69 17747 407 17781
rect -69 17489 407 17523
rect -69 17331 407 17365
rect -69 17073 407 17107
rect -69 16915 407 16949
rect -69 16657 407 16691
rect -69 16499 407 16533
rect -69 16241 407 16275
rect -69 16083 407 16117
rect -69 15825 407 15859
rect 8 14125 42 14601
rect 266 14125 300 14601
rect 424 14125 458 14601
rect 682 14125 716 14601
rect 840 14125 874 14601
rect 1098 14125 1132 14601
rect 1256 14125 1290 14601
rect 1514 14125 1548 14601
rect 1672 14125 1706 14601
rect 1930 14125 1964 14601
rect 2088 14125 2122 14601
rect 2346 14125 2380 14601
rect 613 13541 647 13717
rect 1671 13541 1705 13717
rect 5845 18179 5879 19255
rect 6063 18179 6097 19255
rect 6245 18179 6279 19255
rect 6463 18179 6497 19255
rect 6645 18179 6679 19255
rect 6863 18179 6897 19255
rect 7045 18179 7079 19255
rect 7263 18179 7297 19255
rect 7445 18179 7479 19255
rect 7663 18179 7697 19255
rect 7845 18179 7879 19255
rect 8063 18179 8097 19255
rect 8245 18179 8279 19255
rect 8463 18179 8497 19255
rect 8645 18179 8679 19255
rect 8863 18179 8897 19255
rect 9045 18179 9079 19255
rect 9263 18179 9297 19255
rect 9445 18179 9479 19255
rect 9663 18179 9697 19255
rect 9845 18179 9879 19255
rect 10063 18179 10097 19255
rect 10245 18179 10279 19255
rect 10463 18179 10497 19255
rect 10645 18179 10679 19255
rect 10863 18179 10897 19255
rect 11045 18179 11079 19255
rect 11263 18179 11297 19255
rect 11445 18179 11479 19255
rect 11663 18179 11697 19255
rect 11845 18179 11879 19255
rect 12063 18179 12097 19255
rect 5724 16479 5758 17555
rect 5942 16479 5976 17555
rect 6124 16479 6158 17555
rect 6342 16479 6376 17555
rect 6524 16479 6558 17555
rect 6742 16479 6776 17555
rect 6924 16479 6958 17555
rect 7142 16479 7176 17555
rect 7324 16479 7358 17555
rect 7542 16479 7576 17555
rect 7724 16479 7758 17555
rect 7942 16479 7976 17555
rect 8124 16479 8158 17555
rect 8342 16479 8376 17555
rect 8524 16479 8558 17555
rect 8742 16479 8776 17555
rect 5942 15487 7018 15521
rect 7418 15443 8494 15477
rect 5942 15269 7018 15303
rect 7418 15305 8494 15339
rect 5942 15127 7018 15161
rect 7418 15145 8494 15179
rect 7418 15007 8494 15041
rect 5942 14909 7018 14943
rect 7388 14863 8464 14897
rect 5942 14767 7018 14801
rect 7388 14605 8464 14639
rect 5942 14549 7018 14583
rect 5942 14407 7018 14441
rect 7388 14439 8464 14473
rect 5942 14189 7018 14223
rect 7388 14181 8464 14215
rect 10523 15443 11599 15477
rect 11999 15487 13075 15521
rect 10523 15305 11599 15339
rect 11999 15269 13075 15303
rect 10523 15145 11599 15179
rect 11999 15127 13075 15161
rect 10523 15007 11599 15041
rect 11999 14909 13075 14943
rect 10553 14863 11629 14897
rect 11999 14767 13075 14801
rect 10553 14605 11629 14639
rect 11999 14549 13075 14583
rect 10553 14439 11629 14473
rect 11999 14407 13075 14441
rect 10553 14181 11629 14215
rect 11999 14189 13075 14223
rect 5942 13821 7018 13855
rect 7418 13777 8494 13811
rect 5942 13603 7018 13637
rect 7418 13639 8494 13673
rect 5942 13461 7018 13495
rect 7418 13479 8494 13513
rect 7418 13341 8494 13375
rect 5942 13243 7018 13277
rect 7388 13197 8464 13231
rect 5942 13101 7018 13135
rect 7388 12939 8464 12973
rect 5942 12883 7018 12917
rect 5942 12741 7018 12775
rect 7388 12773 8464 12807
rect 5942 12523 7018 12557
rect 7388 12515 8464 12549
rect 10523 13777 11599 13811
rect 11999 13821 13075 13855
rect 10523 13639 11599 13673
rect 11999 13603 13075 13637
rect 10523 13479 11599 13513
rect 11999 13461 13075 13495
rect 10523 13341 11599 13375
rect 11999 13243 13075 13277
rect 10553 13197 11629 13231
rect 11999 13101 13075 13135
rect 10553 12939 11629 12973
rect 11999 12883 13075 12917
rect 10553 12773 11629 12807
rect 11999 12741 13075 12775
rect 10553 12515 11629 12549
rect 11999 12523 13075 12557
rect 5942 12155 7018 12189
rect 7418 12111 8494 12145
rect 5942 11937 7018 11971
rect 7418 11973 8494 12007
rect 5942 11795 7018 11829
rect 7418 11813 8494 11847
rect 7418 11675 8494 11709
rect 5942 11577 7018 11611
rect 7388 11531 8464 11565
rect 5942 11435 7018 11469
rect 7388 11273 8464 11307
rect 5942 11217 7018 11251
rect 5942 11075 7018 11109
rect 7388 11107 8464 11141
rect 5942 10857 7018 10891
rect 7388 10849 8464 10883
rect 10523 12111 11599 12145
rect 11999 12155 13075 12189
rect 10523 11973 11599 12007
rect 11999 11937 13075 11971
rect 10523 11813 11599 11847
rect 11999 11795 13075 11829
rect 10523 11675 11599 11709
rect 11999 11577 13075 11611
rect 10553 11531 11629 11565
rect 11999 11435 13075 11469
rect 10553 11273 11629 11307
rect 11999 11217 13075 11251
rect 10553 11107 11629 11141
rect 11999 11075 13075 11109
rect 10553 10849 11629 10883
rect 11999 10857 13075 10891
rect 5942 10489 7018 10523
rect 7418 10445 8494 10479
rect 5942 10271 7018 10305
rect 7418 10307 8494 10341
rect 5942 10129 7018 10163
rect 7418 10147 8494 10181
rect 7418 10009 8494 10043
rect 5942 9911 7018 9945
rect 7388 9865 8464 9899
rect 5942 9769 7018 9803
rect 7388 9607 8464 9641
rect 5942 9551 7018 9585
rect 5942 9409 7018 9443
rect 7388 9441 8464 9475
rect 5942 9191 7018 9225
rect 7388 9183 8464 9217
rect 10523 10445 11599 10479
rect 11999 10489 13075 10523
rect 10523 10307 11599 10341
rect 11999 10271 13075 10305
rect 10523 10147 11599 10181
rect 11999 10129 13075 10163
rect 10523 10009 11599 10043
rect 11999 9911 13075 9945
rect 10553 9865 11629 9899
rect 11999 9769 13075 9803
rect 10553 9607 11629 9641
rect 11999 9551 13075 9585
rect 10553 9441 11629 9475
rect 11999 9409 13075 9443
rect 10553 9183 11629 9217
rect 11999 9191 13075 9225
rect 5942 8823 7018 8857
rect 7418 8779 8494 8813
rect 5942 8605 7018 8639
rect 7418 8641 8494 8675
rect 5942 8463 7018 8497
rect 7418 8481 8494 8515
rect 7418 8343 8494 8377
rect 5942 8245 7018 8279
rect 7388 8199 8464 8233
rect 5942 8103 7018 8137
rect 7388 7941 8464 7975
rect 5942 7885 7018 7919
rect 5942 7743 7018 7777
rect 7388 7775 8464 7809
rect 5942 7525 7018 7559
rect 7388 7517 8464 7551
rect 10523 8779 11599 8813
rect 11999 8823 13075 8857
rect 10523 8641 11599 8675
rect 11999 8605 13075 8639
rect 10523 8481 11599 8515
rect 11999 8463 13075 8497
rect 10523 8343 11599 8377
rect 11999 8245 13075 8279
rect 10553 8199 11629 8233
rect 11999 8103 13075 8137
rect 10553 7941 11629 7975
rect 11999 7885 13075 7919
rect 10553 7775 11629 7809
rect 11999 7743 13075 7777
rect 10553 7517 11629 7551
rect 11999 7525 13075 7559
rect 16250 17462 17426 17496
rect 16250 17226 17426 17260
rect 16250 17092 17426 17126
rect 16250 16856 17426 16890
rect 16486 16324 16520 16644
rect 17164 16324 17198 16644
rect 17374 16432 17408 16572
rect 17642 16432 17676 16572
rect 14502 10648 14536 11662
rect 14846 10648 14880 11662
rect 14502 9392 14536 10406
rect 14846 9392 14880 10406
rect 14476 7590 14510 8586
rect 14666 7590 14700 8586
rect 14876 7590 14910 8586
rect 15066 7590 15100 8586
rect 15276 7590 15310 8586
rect 15466 7590 15500 8586
rect 15676 7590 15710 8586
rect 15866 7590 15900 8586
rect 16076 7590 16110 8586
rect 16266 7590 16300 8586
rect 16476 7590 16510 8586
rect 16666 7590 16700 8586
rect 16876 7590 16910 8586
rect 17066 7590 17100 8586
rect 17276 7590 17310 8586
rect 17466 7590 17500 8586
rect 17676 7590 17710 8586
rect 17866 7590 17900 8586
rect 18076 7590 18110 8586
rect 18266 7590 18300 8586
<< pdiffc >>
rect 1340 19110 1374 19186
rect 1798 19110 1832 19186
rect 2040 19110 2074 19186
rect 2498 19110 2532 19186
rect 1340 18326 1374 18802
rect 1798 18326 1832 18802
rect 2040 18326 2074 18802
rect 2498 18326 2532 18802
rect 1340 17542 1374 18018
rect 1798 17542 1832 18018
rect 2040 17542 2074 18018
rect 2498 17542 2532 18018
rect 1340 16758 1374 17234
rect 1798 16758 1832 17234
rect 2040 16758 2074 17234
rect 2498 16758 2532 17234
rect 1340 15974 1374 16450
rect 1798 15974 1832 16450
rect 2040 15974 2074 16450
rect 2498 15974 2532 16450
rect 1340 15590 1374 15666
rect 1798 15590 1832 15666
rect 2040 15590 2074 15666
rect 2498 15590 2532 15666
rect -151 12692 225 12726
rect 485 12692 861 12726
rect 1121 12692 1497 12726
rect 1757 12692 2133 12726
rect -151 12534 225 12568
rect 485 12534 861 12568
rect 1121 12534 1497 12568
rect 1757 12534 2133 12568
rect 733 11735 767 11887
rect 2185 11735 2219 11887
rect 355 10323 389 10985
rect 967 10323 1001 10985
rect 1349 10903 1383 10979
rect 2207 10903 2241 10979
rect 1275 10137 1309 10587
rect 2209 10137 2243 10587
rect 1109 8764 1143 9240
rect 1567 8764 1601 9240
rect 1809 8764 1843 9240
rect 2267 8764 2301 9240
rect 1109 7980 1143 8456
rect 1567 7980 1601 8456
rect 1809 7980 1843 8456
rect 2267 7980 2301 8456
rect 3036 19126 3070 19202
rect 3494 19126 3528 19202
rect 3736 19126 3770 19202
rect 4194 19126 4228 19202
rect 3036 18342 3070 18818
rect 3494 18342 3528 18818
rect 3736 18342 3770 18818
rect 4194 18342 4228 18818
rect 3036 17558 3070 18034
rect 3494 17558 3528 18034
rect 3736 17558 3770 18034
rect 4194 17558 4228 18034
rect 3036 16774 3070 17250
rect 3494 16774 3528 17250
rect 3736 16774 3770 17250
rect 4194 16774 4228 17250
rect 3036 15990 3070 16466
rect 3494 15990 3528 16466
rect 3736 15990 3770 16466
rect 4194 15990 4228 16466
rect 3036 15206 3070 15682
rect 3494 15206 3528 15682
rect 3736 15206 3770 15682
rect 4194 15206 4228 15682
rect 3036 14422 3070 14898
rect 3494 14422 3528 14898
rect 3736 14422 3770 14898
rect 4194 14422 4228 14898
rect 3036 13638 3070 14114
rect 3494 13638 3528 14114
rect 3736 13638 3770 14114
rect 4194 13638 4228 14114
rect 3036 12854 3070 13330
rect 3494 12854 3528 13330
rect 3736 12854 3770 13330
rect 4194 12854 4228 13330
rect 3036 12070 3070 12546
rect 3494 12070 3528 12546
rect 3736 12070 3770 12546
rect 4194 12070 4228 12546
rect 3036 11286 3070 11762
rect 3494 11286 3528 11762
rect 3736 11286 3770 11762
rect 4194 11286 4228 11762
rect 3036 10502 3070 10978
rect 3494 10502 3528 10978
rect 3736 10502 3770 10978
rect 4194 10502 4228 10978
rect 3036 9718 3070 10194
rect 3494 9718 3528 10194
rect 3736 9718 3770 10194
rect 4194 9718 4228 10194
rect 3036 8934 3070 9410
rect 3494 8934 3528 9410
rect 3736 8934 3770 9410
rect 4194 8934 4228 9410
rect 3036 8150 3070 8626
rect 3494 8150 3528 8626
rect 3736 8150 3770 8626
rect 4194 8150 4228 8626
rect 3036 7766 3070 7842
rect 3494 7766 3528 7842
rect 3736 7766 3770 7842
rect 4194 7766 4228 7842
rect 9368 17126 9402 17302
rect 9586 17126 9620 17302
rect 9768 17126 9802 17302
rect 9986 17126 10020 17302
rect 10627 17097 10661 17273
rect 10845 17097 10879 17273
rect 11027 17097 11061 17273
rect 11245 17097 11279 17273
rect 11427 17097 11461 17273
rect 11645 17097 11679 17273
rect 11827 17097 11861 17273
rect 12045 17097 12079 17273
rect 9075 15518 9251 15552
rect 9075 15300 9251 15334
rect 9075 15110 9251 15144
rect 9075 14892 9251 14926
rect 9075 14664 9251 14698
rect 9075 14206 9251 14240
rect 9766 15518 9942 15552
rect 9766 15300 9942 15334
rect 9766 15110 9942 15144
rect 9766 14892 9942 14926
rect 9766 14664 9942 14698
rect 9766 14206 9942 14240
rect 9075 13852 9251 13886
rect 9075 13634 9251 13668
rect 9075 13444 9251 13478
rect 9075 13226 9251 13260
rect 9075 12998 9251 13032
rect 9075 12540 9251 12574
rect 9766 13852 9942 13886
rect 9766 13634 9942 13668
rect 9766 13444 9942 13478
rect 9766 13226 9942 13260
rect 9766 12998 9942 13032
rect 9766 12540 9942 12574
rect 9075 12186 9251 12220
rect 9075 11968 9251 12002
rect 9075 11778 9251 11812
rect 9075 11560 9251 11594
rect 9075 11332 9251 11366
rect 9075 10874 9251 10908
rect 9766 12186 9942 12220
rect 9766 11968 9942 12002
rect 9766 11778 9942 11812
rect 9766 11560 9942 11594
rect 9766 11332 9942 11366
rect 9766 10874 9942 10908
rect 9075 10520 9251 10554
rect 9075 10302 9251 10336
rect 9075 10112 9251 10146
rect 9075 9894 9251 9928
rect 9075 9666 9251 9700
rect 9075 9208 9251 9242
rect 9766 10520 9942 10554
rect 9766 10302 9942 10336
rect 9766 10112 9942 10146
rect 9766 9894 9942 9928
rect 9766 9666 9942 9700
rect 9766 9208 9942 9242
rect 9075 8854 9251 8888
rect 9075 8636 9251 8670
rect 9075 8446 9251 8480
rect 9075 8228 9251 8262
rect 9075 8000 9251 8034
rect 9075 7542 9251 7576
rect 9766 8854 9942 8888
rect 9766 8636 9942 8670
rect 9766 8446 9942 8480
rect 9766 8228 9942 8262
rect 9766 8000 9942 8034
rect 9766 7542 9942 7576
rect 15055 15977 15089 17673
rect 15183 15977 15217 17673
rect 14994 13468 15148 13502
rect 15494 13468 15648 13502
rect 15994 13468 16148 13502
rect 16494 13468 16648 13502
rect 16994 13468 17148 13502
rect 17494 13468 17648 13502
rect 14994 12632 15148 12666
rect 15494 12632 15648 12666
rect 15994 12632 16148 12666
rect 16494 12632 16648 12666
rect 16994 12632 17148 12666
rect 17494 12632 17648 12666
rect 17098 11313 18108 11347
rect 17098 11181 18108 11215
rect 17041 10246 18231 10280
rect 17041 9934 18231 9968
rect 17041 9646 18231 9680
rect 17041 9334 18231 9368
<< psubdiff >>
rect 5460 19716 5590 19740
rect -588 19530 -564 19683
rect 4357 19613 4673 19683
rect 4357 19530 4507 19613
rect -560 19401 -436 19530
rect -269 19110 -99 19198
rect 576 19110 633 19198
rect -269 19100 -200 19110
rect 582 19035 633 19110
rect 582 15702 633 15793
rect -200 15674 -115 15702
rect -269 15614 -115 15674
rect 560 15614 633 15702
rect -203 14773 -4 14846
rect 2394 14773 2549 14846
rect -203 14754 -115 14773
rect 2461 14770 2549 14773
rect -203 13903 -115 14079
rect 2461 14007 2549 14095
rect 2461 13905 2551 14007
rect 1804 13903 1897 13905
rect -237 13809 -213 13903
rect 393 13869 595 13903
rect 1723 13869 1897 13903
rect 393 13809 533 13869
rect 1785 13829 1897 13869
rect 2527 13829 2551 13905
rect 499 13807 533 13809
rect 1785 13807 1819 13829
rect 499 13389 533 13451
rect 1785 13389 1819 13451
rect 499 13355 595 13389
rect 1723 13355 1819 13389
rect 2467 12860 2584 12884
rect 290 12179 314 12294
rect 2111 12179 2467 12294
rect 2467 9748 2584 9772
rect -560 7379 -436 7535
rect -561 7226 -537 7379
rect 4384 7324 4507 7379
rect 12542 19716 12672 19740
rect 5590 19565 5662 19689
rect 12451 19565 12542 19689
rect 5590 16142 5655 16266
rect 12444 16142 12542 16266
rect 5460 16118 5590 16142
rect 12542 16118 12672 16142
rect 14352 18214 18330 18222
rect 14352 18198 14644 18214
rect 8549 15840 10468 15931
rect 8549 15720 8672 15840
rect 4384 7226 4673 7324
rect 5452 15692 5734 15720
rect 5606 15630 5734 15692
rect 8648 15630 8672 15720
rect 10345 15720 10468 15840
rect 8549 15625 8672 15630
rect 8641 14289 8759 14313
rect 8641 14147 8759 14171
rect 10345 15630 10369 15720
rect 13283 15692 13565 15720
rect 13283 15630 13411 15692
rect 10345 15625 10468 15630
rect 10258 14289 10376 14313
rect 10258 14147 10376 14171
rect 5606 13964 5734 14054
rect 8648 13964 8672 14054
rect 8641 12623 8759 12647
rect 8641 12481 8759 12505
rect 10345 13964 10369 14054
rect 13283 13964 13411 14054
rect 10258 12623 10376 12647
rect 10258 12481 10376 12505
rect 5606 12298 5734 12388
rect 8648 12298 8672 12388
rect 8641 10957 8759 10981
rect 8641 10815 8759 10839
rect 10345 12298 10369 12388
rect 13283 12298 13411 12388
rect 10258 10957 10376 10981
rect 10258 10815 10376 10839
rect 5606 10632 5734 10722
rect 8648 10632 8672 10722
rect 8641 9291 8759 9315
rect 8641 9149 8759 9173
rect 10345 10632 10369 10722
rect 13283 10632 13411 10722
rect 10258 9291 10376 9315
rect 10258 9149 10376 9173
rect 5606 8966 5734 9056
rect 8648 8966 8672 9056
rect 8641 7625 8759 7649
rect 8641 7483 8759 7507
rect 10345 8966 10369 9056
rect 13283 8966 13411 9056
rect 10258 7625 10376 7649
rect 10258 7483 10376 7507
rect 5606 7284 5735 7292
rect 5452 7212 5735 7284
rect 13377 7284 13411 7292
rect 14530 18057 14644 18198
rect 18041 18198 18330 18214
rect 18041 18057 18152 18198
rect 15808 17618 15928 17658
rect 15882 17590 15928 17618
rect 17742 17618 17896 17658
rect 17742 17590 17822 17618
rect 15882 16052 15954 16092
rect 15808 16024 15954 16052
rect 17648 16024 17724 16092
rect 17768 16052 17822 16092
rect 17768 16024 17896 16052
rect 14530 15597 18152 15605
rect 14530 15473 14634 15597
rect 14352 15440 14634 15473
rect 18031 15473 18152 15597
rect 18031 15440 18330 15473
rect 14387 13772 14444 13864
rect 18497 13772 18637 13864
rect 14387 13722 14466 13772
rect 18551 13756 18637 13772
rect 14387 11848 14466 12335
rect 14387 11843 14484 11848
rect 14388 11814 14484 11843
rect 14898 11814 14994 11848
rect 14388 11752 14422 11814
rect 14960 11752 14994 11814
rect 14388 9240 14422 9302
rect 14960 9240 14994 9302
rect 14388 9206 14484 9240
rect 14898 9206 14994 9240
rect 14424 8850 14558 9206
rect 14298 8766 14383 8850
rect 18441 8766 18551 8850
rect 14298 8693 14380 8766
rect 18404 8675 18551 8766
rect 14298 7430 14380 7529
rect 18486 7511 18551 8675
rect 18404 7430 18551 7511
rect 14298 7346 14383 7430
rect 18441 7350 18551 7430
rect 18441 7346 18637 7350
rect 18464 7326 18637 7346
rect 13377 7212 13565 7284
<< nsubdiff >>
rect 1057 19363 1117 19397
rect 2631 19363 2691 19397
rect 1057 19337 1091 19363
rect 2657 19337 2691 19363
rect 1057 15427 1091 15453
rect 2657 15427 2691 15453
rect 1057 15393 1117 15427
rect 2631 15393 2691 15427
rect 2883 19379 2943 19413
rect 4314 19379 4374 19413
rect 2883 19353 2917 19379
rect -346 12806 -250 12840
rect 2232 12806 2328 12840
rect -346 12744 -312 12806
rect 2294 12744 2328 12806
rect -346 12454 -312 12516
rect 2294 12454 2328 12516
rect -346 12420 -250 12454
rect 2232 12420 2328 12454
rect 619 12048 715 12082
rect 2237 12048 2333 12082
rect 619 11986 653 12048
rect 2299 11986 2333 12048
rect 619 11574 653 11636
rect 2299 11574 2333 11636
rect 619 11540 715 11574
rect 2237 11540 2333 11574
rect 241 11170 301 11204
rect 2297 11170 2357 11204
rect 241 11144 275 11170
rect 2323 11144 2357 11170
rect 241 9943 275 9969
rect 2323 9943 2357 9969
rect 241 9909 301 9943
rect 2297 9909 2357 9943
rect 973 9391 1033 9425
rect 2373 9391 2433 9425
rect 973 9365 1007 9391
rect 2399 9365 2433 9391
rect 973 7817 1007 7843
rect 2399 7817 2433 7843
rect 973 7783 1033 7817
rect 2373 7783 2433 7817
rect 4340 19353 4374 19379
rect 2883 7612 2917 7638
rect 4340 7612 4374 7638
rect 2883 7578 2943 7612
rect 4314 7578 4374 7612
rect 9108 17585 9168 17619
rect 10222 17585 10282 17619
rect 9108 17559 9142 17585
rect 10248 17559 10282 17585
rect 9108 16837 9142 16863
rect 10248 16837 10282 16863
rect 9108 16803 9168 16837
rect 10222 16803 10282 16837
rect 10401 17574 10461 17608
rect 12244 17574 12304 17608
rect 10401 17548 10435 17574
rect 12270 17548 12304 17574
rect 10401 16757 10435 16783
rect 12270 16757 12304 16783
rect 10401 16723 10461 16757
rect 12244 16723 12304 16757
rect 8861 15652 8921 15686
rect 9407 15652 9467 15686
rect 8861 15626 8895 15652
rect 9433 15626 9467 15652
rect 8861 14126 8895 14152
rect 9433 14126 9467 14152
rect 8861 14092 8921 14126
rect 9407 14092 9467 14126
rect 9550 15652 9610 15686
rect 10096 15652 10156 15686
rect 9550 15626 9584 15652
rect 10122 15626 10156 15652
rect 9550 14126 9584 14152
rect 10122 14126 10156 14152
rect 9550 14092 9610 14126
rect 10096 14092 10156 14126
rect 8861 13986 8921 14020
rect 9407 13986 9467 14020
rect 8861 13960 8895 13986
rect 9433 13960 9467 13986
rect 8861 12460 8895 12486
rect 9433 12460 9467 12486
rect 8861 12426 8921 12460
rect 9407 12426 9467 12460
rect 9550 13986 9610 14020
rect 10096 13986 10156 14020
rect 9550 13960 9584 13986
rect 10122 13960 10156 13986
rect 9550 12460 9584 12486
rect 10122 12460 10156 12486
rect 9550 12426 9610 12460
rect 10096 12426 10156 12460
rect 8861 12320 8921 12354
rect 9407 12320 9467 12354
rect 8861 12294 8895 12320
rect 9433 12294 9467 12320
rect 8861 10794 8895 10820
rect 9433 10794 9467 10820
rect 8861 10760 8921 10794
rect 9407 10760 9467 10794
rect 9550 12320 9610 12354
rect 10096 12320 10156 12354
rect 9550 12294 9584 12320
rect 10122 12294 10156 12320
rect 9550 10794 9584 10820
rect 10122 10794 10156 10820
rect 9550 10760 9610 10794
rect 10096 10760 10156 10794
rect 8861 10654 8921 10688
rect 9407 10654 9467 10688
rect 8861 10628 8895 10654
rect 9433 10628 9467 10654
rect 8861 9128 8895 9154
rect 9433 9128 9467 9154
rect 8861 9094 8921 9128
rect 9407 9094 9467 9128
rect 9550 10654 9610 10688
rect 10096 10654 10156 10688
rect 9550 10628 9584 10654
rect 10122 10628 10156 10654
rect 9550 9128 9584 9154
rect 10122 9128 10156 9154
rect 9550 9094 9610 9128
rect 10096 9094 10156 9128
rect 8861 8988 8921 9022
rect 9407 8988 9467 9022
rect 8861 8962 8895 8988
rect 9433 8962 9467 8988
rect 8861 7462 8895 7488
rect 9433 7462 9467 7488
rect 8861 7428 8921 7462
rect 9407 7428 9467 7462
rect 9550 8988 9610 9022
rect 10096 8988 10156 9022
rect 9550 8962 9584 8988
rect 10122 8962 10156 8988
rect 9550 7462 9584 7488
rect 10122 7462 10156 7488
rect 9550 7428 9610 7462
rect 10096 7428 10156 7462
rect 14750 17836 14810 17870
rect 15463 17836 15523 17870
rect 14750 17810 14784 17836
rect 15489 17810 15523 17836
rect 14750 15823 14784 15849
rect 15489 15823 15523 15849
rect 14750 15789 14810 15823
rect 15463 15789 15523 15823
rect 14764 13644 14824 13678
rect 17845 13644 17905 13678
rect 14764 13618 14798 13644
rect 17871 13618 17905 13644
rect 14764 12491 14798 12517
rect 17871 12491 17905 12517
rect 14764 12457 14824 12491
rect 17845 12457 17905 12491
rect 16903 11427 16999 11461
rect 18207 11427 18303 11461
rect 16903 11365 16937 11427
rect 18269 11365 18303 11427
rect 16903 11101 16937 11163
rect 18269 11101 18303 11163
rect 16903 11067 16999 11101
rect 18207 11067 18303 11101
rect 16843 10407 16903 10441
rect 18382 10407 18442 10441
rect 16843 10381 16877 10407
rect 18408 10381 18442 10407
rect 16843 9203 16877 9229
rect 18408 9203 18442 9229
rect 16843 9169 16903 9203
rect 18382 9169 18442 9203
<< psubdiffcont >>
rect -564 19530 4357 19683
rect -560 7535 -436 19401
rect -99 19110 576 19198
rect -269 15674 -200 19100
rect 582 15793 633 19035
rect -115 15614 560 15702
rect -4 14773 2394 14846
rect -203 14079 -115 14754
rect 2461 14095 2549 14770
rect -213 13809 393 13903
rect 595 13869 1723 13903
rect 1897 13829 2527 13905
rect 499 13451 533 13807
rect 1785 13451 1819 13807
rect 595 13355 1723 13389
rect 314 12179 2111 12294
rect 2467 9772 2584 12860
rect -537 7226 4384 7379
rect 4507 7324 4673 19613
rect 5460 16142 5590 19716
rect 5662 19565 12451 19689
rect 5655 16142 12444 16266
rect 12542 16142 12672 19716
rect 5452 7284 5606 15692
rect 5734 15630 8648 15720
rect 8641 14171 8759 14289
rect 10369 15630 13283 15720
rect 10258 14171 10376 14289
rect 5734 13964 8648 14054
rect 8641 12505 8759 12623
rect 10369 13964 13283 14054
rect 10258 12505 10376 12623
rect 5734 12298 8648 12388
rect 8641 10839 8759 10957
rect 10369 12298 13283 12388
rect 10258 10839 10376 10957
rect 5734 10632 8648 10722
rect 8641 9173 8759 9291
rect 10369 10632 13283 10722
rect 10258 9173 10376 9291
rect 5734 8966 8648 9056
rect 8641 7507 8759 7625
rect 10369 8966 13283 9056
rect 10258 7507 10376 7625
rect 5735 7212 13377 7292
rect 13411 7284 13565 15692
rect 14352 15473 14530 18198
rect 14644 18057 18041 18214
rect 15808 16052 15882 17618
rect 15928 17590 17742 17658
rect 15954 16024 17648 16092
rect 17724 16024 17768 16092
rect 17822 16052 17896 17618
rect 14634 15440 18031 15597
rect 18152 15473 18330 18198
rect 14444 13772 18497 13864
rect 14387 12335 14466 13722
rect 14484 11814 14898 11848
rect 14388 9302 14422 11752
rect 14960 9302 14994 11752
rect 14484 9206 14898 9240
rect 14383 8766 18441 8850
rect 14298 7529 14380 8693
rect 18404 7511 18486 8675
rect 14383 7346 18441 7430
rect 18551 7350 18637 13756
<< nsubdiffcont >>
rect 1117 19363 2631 19397
rect 1057 15453 1091 19337
rect 2657 15453 2691 19337
rect 1117 15393 2631 15427
rect 2943 19379 4314 19413
rect -250 12806 2232 12840
rect -346 12516 -312 12744
rect 2294 12516 2328 12744
rect -250 12420 2232 12454
rect 715 12048 2237 12082
rect 619 11636 653 11986
rect 2299 11636 2333 11986
rect 715 11540 2237 11574
rect 301 11170 2297 11204
rect 241 9969 275 11144
rect 2323 9969 2357 11144
rect 301 9909 2297 9943
rect 1033 9391 2373 9425
rect 973 7843 1007 9365
rect 2399 7843 2433 9365
rect 1033 7783 2373 7817
rect 2883 7638 2917 19353
rect 4340 7638 4374 19353
rect 2943 7578 4314 7612
rect 9168 17585 10222 17619
rect 9108 16863 9142 17559
rect 10248 16863 10282 17559
rect 9168 16803 10222 16837
rect 10461 17574 12244 17608
rect 10401 16783 10435 17548
rect 12270 16783 12304 17548
rect 10461 16723 12244 16757
rect 8921 15652 9407 15686
rect 8861 14152 8895 15626
rect 9433 14152 9467 15626
rect 8921 14092 9407 14126
rect 9610 15652 10096 15686
rect 9550 14152 9584 15626
rect 10122 14152 10156 15626
rect 9610 14092 10096 14126
rect 8921 13986 9407 14020
rect 8861 12486 8895 13960
rect 9433 12486 9467 13960
rect 8921 12426 9407 12460
rect 9610 13986 10096 14020
rect 9550 12486 9584 13960
rect 10122 12486 10156 13960
rect 9610 12426 10096 12460
rect 8921 12320 9407 12354
rect 8861 10820 8895 12294
rect 9433 10820 9467 12294
rect 8921 10760 9407 10794
rect 9610 12320 10096 12354
rect 9550 10820 9584 12294
rect 10122 10820 10156 12294
rect 9610 10760 10096 10794
rect 8921 10654 9407 10688
rect 8861 9154 8895 10628
rect 9433 9154 9467 10628
rect 8921 9094 9407 9128
rect 9610 10654 10096 10688
rect 9550 9154 9584 10628
rect 10122 9154 10156 10628
rect 9610 9094 10096 9128
rect 8921 8988 9407 9022
rect 8861 7488 8895 8962
rect 9433 7488 9467 8962
rect 8921 7428 9407 7462
rect 9610 8988 10096 9022
rect 9550 7488 9584 8962
rect 10122 7488 10156 8962
rect 9610 7428 10096 7462
rect 14810 17836 15463 17870
rect 14750 15849 14784 17810
rect 15489 15849 15523 17810
rect 14810 15789 15463 15823
rect 14824 13644 17845 13678
rect 14764 12517 14798 13618
rect 17871 12517 17905 13618
rect 14824 12457 17845 12491
rect 16999 11427 18207 11461
rect 16903 11163 16937 11365
rect 18269 11163 18303 11365
rect 16999 11067 18207 11101
rect 16903 10407 18382 10441
rect 16843 9229 16877 10381
rect 18408 9229 18442 10381
rect 16903 9169 18382 9203
<< poly >>
rect -169 18967 -81 18983
rect -169 18799 -153 18967
rect -119 18799 -81 18967
rect -169 18783 -81 18799
rect 419 18967 507 18983
rect 419 18799 457 18967
rect 491 18799 507 18967
rect 419 18783 507 18799
rect -169 18551 -81 18567
rect -169 18383 -153 18551
rect -119 18383 -81 18551
rect -169 18367 -81 18383
rect 419 18551 507 18567
rect 419 18383 457 18551
rect 491 18383 507 18551
rect 419 18367 507 18383
rect -169 18135 -81 18151
rect -169 17967 -153 18135
rect -119 17967 -81 18135
rect -169 17951 -81 17967
rect 419 18135 507 18151
rect 419 17967 457 18135
rect 491 17967 507 18135
rect 419 17951 507 17967
rect -169 17719 -81 17735
rect -169 17551 -153 17719
rect -119 17551 -81 17719
rect -169 17535 -81 17551
rect 419 17719 507 17735
rect 419 17551 457 17719
rect 491 17551 507 17719
rect 419 17535 507 17551
rect -169 17303 -81 17319
rect -169 17135 -153 17303
rect -119 17135 -81 17303
rect -169 17119 -81 17135
rect 419 17303 507 17319
rect 419 17135 457 17303
rect 491 17135 507 17303
rect 419 17119 507 17135
rect -169 16887 -81 16903
rect -169 16719 -153 16887
rect -119 16719 -81 16887
rect -169 16703 -81 16719
rect 419 16887 507 16903
rect 419 16719 457 16887
rect 491 16719 507 16887
rect 419 16703 507 16719
rect -169 16471 -81 16487
rect -169 16303 -153 16471
rect -119 16303 -81 16471
rect -169 16287 -81 16303
rect 419 16471 507 16487
rect 419 16303 457 16471
rect 491 16303 507 16471
rect 419 16287 507 16303
rect -169 16055 -81 16071
rect -169 15887 -153 16055
rect -119 15887 -81 16055
rect -169 15871 -81 15887
rect 419 16055 507 16071
rect 419 15887 457 16055
rect 491 15887 507 16055
rect 419 15871 507 15887
rect 1386 19279 1786 19295
rect 1386 19245 1402 19279
rect 1770 19245 1786 19279
rect 1386 19198 1786 19245
rect 2086 19279 2486 19295
rect 2086 19245 2102 19279
rect 2470 19245 2486 19279
rect 2086 19198 2486 19245
rect 1386 19051 1786 19098
rect 1386 19017 1402 19051
rect 1770 19017 1786 19051
rect 1386 19001 1786 19017
rect 2086 19051 2486 19098
rect 2086 19017 2102 19051
rect 2470 19017 2486 19051
rect 2086 19001 2486 19017
rect 1386 18895 1786 18911
rect 1386 18861 1402 18895
rect 1770 18861 1786 18895
rect 1386 18814 1786 18861
rect 2086 18895 2486 18911
rect 2086 18861 2102 18895
rect 2470 18861 2486 18895
rect 2086 18814 2486 18861
rect 1386 18267 1786 18314
rect 1386 18233 1402 18267
rect 1770 18233 1786 18267
rect 1386 18217 1786 18233
rect 2086 18267 2486 18314
rect 2086 18233 2102 18267
rect 2470 18233 2486 18267
rect 2086 18217 2486 18233
rect 1386 18111 1786 18127
rect 1386 18077 1402 18111
rect 1770 18077 1786 18111
rect 1386 18030 1786 18077
rect 2086 18111 2486 18127
rect 2086 18077 2102 18111
rect 2470 18077 2486 18111
rect 2086 18030 2486 18077
rect 1386 17483 1786 17530
rect 1386 17449 1402 17483
rect 1770 17449 1786 17483
rect 1386 17433 1786 17449
rect 2086 17483 2486 17530
rect 2086 17449 2102 17483
rect 2470 17449 2486 17483
rect 2086 17433 2486 17449
rect 1386 17327 1786 17343
rect 1386 17293 1402 17327
rect 1770 17293 1786 17327
rect 1386 17246 1786 17293
rect 2086 17327 2486 17343
rect 2086 17293 2102 17327
rect 2470 17293 2486 17327
rect 2086 17246 2486 17293
rect 1386 16699 1786 16746
rect 1386 16665 1402 16699
rect 1770 16665 1786 16699
rect 1386 16649 1786 16665
rect 2086 16699 2486 16746
rect 2086 16665 2102 16699
rect 2470 16665 2486 16699
rect 2086 16649 2486 16665
rect 1386 16543 1786 16559
rect 1386 16509 1402 16543
rect 1770 16509 1786 16543
rect 1386 16462 1786 16509
rect 2086 16543 2486 16559
rect 2086 16509 2102 16543
rect 2470 16509 2486 16543
rect 2086 16462 2486 16509
rect 1386 15915 1786 15962
rect 1386 15881 1402 15915
rect 1770 15881 1786 15915
rect 1386 15865 1786 15881
rect 2086 15915 2486 15962
rect 2086 15881 2102 15915
rect 2470 15881 2486 15915
rect 2086 15865 2486 15881
rect 1386 15759 1786 15775
rect 1386 15725 1402 15759
rect 1770 15725 1786 15759
rect 1386 15678 1786 15725
rect 2086 15759 2486 15775
rect 2086 15725 2102 15759
rect 2470 15725 2486 15759
rect 2086 15678 2486 15725
rect 1386 15531 1786 15578
rect 1386 15497 1402 15531
rect 1770 15497 1786 15531
rect 1386 15481 1786 15497
rect 2086 15531 2486 15578
rect 2086 15497 2102 15531
rect 2470 15497 2486 15531
rect 2086 15481 2486 15497
rect 54 14685 254 14701
rect 54 14651 70 14685
rect 238 14651 254 14685
rect 54 14613 254 14651
rect 470 14685 670 14701
rect 470 14651 486 14685
rect 654 14651 670 14685
rect 470 14613 670 14651
rect 886 14685 1086 14701
rect 886 14651 902 14685
rect 1070 14651 1086 14685
rect 886 14613 1086 14651
rect 1302 14685 1502 14701
rect 1302 14651 1318 14685
rect 1486 14651 1502 14685
rect 1302 14613 1502 14651
rect 1718 14685 1918 14701
rect 1718 14651 1734 14685
rect 1902 14651 1918 14685
rect 1718 14613 1918 14651
rect 2134 14685 2334 14701
rect 2134 14651 2150 14685
rect 2318 14651 2334 14685
rect 2134 14613 2334 14651
rect 54 14075 254 14113
rect 54 14041 70 14075
rect 238 14041 254 14075
rect 54 14025 254 14041
rect 470 14075 670 14113
rect 470 14041 486 14075
rect 654 14041 670 14075
rect 470 14025 670 14041
rect 886 14075 1086 14113
rect 886 14041 902 14075
rect 1070 14041 1086 14075
rect 886 14025 1086 14041
rect 1302 14075 1502 14113
rect 1302 14041 1318 14075
rect 1486 14041 1502 14075
rect 1302 14025 1502 14041
rect 1718 14075 1918 14113
rect 1718 14041 1734 14075
rect 1902 14041 1918 14075
rect 1718 14025 1918 14041
rect 2134 14075 2334 14113
rect 2134 14041 2150 14075
rect 2318 14041 2334 14075
rect 2134 14025 2334 14041
rect 659 13801 1659 13817
rect 659 13767 675 13801
rect 1643 13767 1659 13801
rect 659 13729 1659 13767
rect 659 13491 1659 13529
rect 659 13457 675 13491
rect 1643 13457 1659 13491
rect 659 13441 1659 13457
rect -260 12664 -163 12680
rect -260 12596 -244 12664
rect -210 12596 -163 12664
rect -260 12580 -163 12596
rect 237 12664 334 12680
rect 237 12596 284 12664
rect 318 12596 334 12664
rect 237 12580 334 12596
rect 376 12664 473 12680
rect 376 12596 392 12664
rect 426 12596 473 12664
rect 376 12580 473 12596
rect 873 12664 970 12680
rect 873 12596 920 12664
rect 954 12596 970 12664
rect 873 12580 970 12596
rect 1012 12664 1109 12680
rect 1012 12596 1028 12664
rect 1062 12596 1109 12664
rect 1012 12580 1109 12596
rect 1509 12664 1606 12680
rect 1509 12596 1556 12664
rect 1590 12596 1606 12664
rect 1509 12580 1606 12596
rect 1648 12664 1745 12680
rect 1648 12596 1664 12664
rect 1698 12596 1745 12664
rect 1648 12580 1745 12596
rect 2145 12664 2242 12680
rect 2145 12596 2192 12664
rect 2226 12596 2242 12664
rect 2145 12580 2242 12596
rect 779 11980 2173 11996
rect 779 11946 795 11980
rect 2157 11946 2173 11980
rect 779 11899 2173 11946
rect 779 11676 2173 11723
rect 779 11642 795 11676
rect 2157 11642 2173 11676
rect 779 11626 2173 11642
rect 401 11078 955 11094
rect 401 11044 417 11078
rect 939 11044 955 11078
rect 401 10997 955 11044
rect 1395 11072 2195 11088
rect 1395 11038 1411 11072
rect 2179 11038 2195 11072
rect 1395 10991 2195 11038
rect 1395 10844 2195 10891
rect 1395 10810 1411 10844
rect 2179 10810 2195 10844
rect 1395 10794 2195 10810
rect 1321 10680 2197 10696
rect 1321 10646 1337 10680
rect 2181 10646 2197 10680
rect 1321 10599 2197 10646
rect 401 10264 955 10311
rect 401 10230 417 10264
rect 939 10230 955 10264
rect 401 10214 955 10230
rect 1321 10078 2197 10125
rect 1321 10044 1337 10078
rect 2181 10044 2197 10078
rect 1321 10028 2197 10044
rect 1155 9333 1555 9349
rect 1155 9299 1171 9333
rect 1539 9299 1555 9333
rect 1155 9252 1555 9299
rect 1855 9333 2255 9349
rect 1855 9299 1871 9333
rect 2239 9299 2255 9333
rect 1855 9252 2255 9299
rect 1155 8705 1555 8752
rect 1155 8671 1171 8705
rect 1539 8671 1555 8705
rect 1155 8655 1555 8671
rect 1855 8705 2255 8752
rect 1855 8671 1871 8705
rect 2239 8671 2255 8705
rect 1855 8655 2255 8671
rect 1155 8549 1555 8565
rect 1155 8515 1171 8549
rect 1539 8515 1555 8549
rect 1155 8468 1555 8515
rect 1855 8549 2255 8565
rect 1855 8515 1871 8549
rect 2239 8515 2255 8549
rect 1855 8468 2255 8515
rect 1155 7921 1555 7968
rect 1155 7887 1171 7921
rect 1539 7887 1555 7921
rect 1155 7871 1555 7887
rect 1855 7921 2255 7968
rect 1855 7887 1871 7921
rect 2239 7887 2255 7921
rect 1855 7871 2255 7887
rect 3082 19295 3482 19311
rect 3082 19261 3098 19295
rect 3466 19261 3482 19295
rect 3082 19214 3482 19261
rect 3782 19295 4182 19311
rect 3782 19261 3798 19295
rect 4166 19261 4182 19295
rect 3782 19214 4182 19261
rect 3082 19067 3482 19114
rect 3082 19033 3098 19067
rect 3466 19033 3482 19067
rect 3082 19017 3482 19033
rect 3782 19067 4182 19114
rect 3782 19033 3798 19067
rect 4166 19033 4182 19067
rect 3782 19017 4182 19033
rect 3082 18911 3482 18927
rect 3082 18877 3098 18911
rect 3466 18877 3482 18911
rect 3082 18830 3482 18877
rect 3782 18911 4182 18927
rect 3782 18877 3798 18911
rect 4166 18877 4182 18911
rect 3782 18830 4182 18877
rect 3082 18283 3482 18330
rect 3082 18249 3098 18283
rect 3466 18249 3482 18283
rect 3082 18233 3482 18249
rect 3782 18283 4182 18330
rect 3782 18249 3798 18283
rect 4166 18249 4182 18283
rect 3782 18233 4182 18249
rect 3082 18127 3482 18143
rect 3082 18093 3098 18127
rect 3466 18093 3482 18127
rect 3082 18046 3482 18093
rect 3782 18127 4182 18143
rect 3782 18093 3798 18127
rect 4166 18093 4182 18127
rect 3782 18046 4182 18093
rect 3082 17499 3482 17546
rect 3082 17465 3098 17499
rect 3466 17465 3482 17499
rect 3082 17449 3482 17465
rect 3782 17499 4182 17546
rect 3782 17465 3798 17499
rect 4166 17465 4182 17499
rect 3782 17449 4182 17465
rect 3082 17343 3482 17359
rect 3082 17309 3098 17343
rect 3466 17309 3482 17343
rect 3082 17262 3482 17309
rect 3782 17343 4182 17359
rect 3782 17309 3798 17343
rect 4166 17309 4182 17343
rect 3782 17262 4182 17309
rect 3082 16715 3482 16762
rect 3082 16681 3098 16715
rect 3466 16681 3482 16715
rect 3082 16665 3482 16681
rect 3782 16715 4182 16762
rect 3782 16681 3798 16715
rect 4166 16681 4182 16715
rect 3782 16665 4182 16681
rect 3082 16559 3482 16575
rect 3082 16525 3098 16559
rect 3466 16525 3482 16559
rect 3082 16478 3482 16525
rect 3782 16559 4182 16575
rect 3782 16525 3798 16559
rect 4166 16525 4182 16559
rect 3782 16478 4182 16525
rect 3082 15931 3482 15978
rect 3082 15897 3098 15931
rect 3466 15897 3482 15931
rect 3082 15881 3482 15897
rect 3782 15931 4182 15978
rect 3782 15897 3798 15931
rect 4166 15897 4182 15931
rect 3782 15881 4182 15897
rect 3082 15775 3482 15791
rect 3082 15741 3098 15775
rect 3466 15741 3482 15775
rect 3082 15694 3482 15741
rect 3782 15775 4182 15791
rect 3782 15741 3798 15775
rect 4166 15741 4182 15775
rect 3782 15694 4182 15741
rect 3082 15147 3482 15194
rect 3082 15113 3098 15147
rect 3466 15113 3482 15147
rect 3082 15097 3482 15113
rect 3782 15147 4182 15194
rect 3782 15113 3798 15147
rect 4166 15113 4182 15147
rect 3782 15097 4182 15113
rect 3082 14991 3482 15007
rect 3082 14957 3098 14991
rect 3466 14957 3482 14991
rect 3082 14910 3482 14957
rect 3782 14991 4182 15007
rect 3782 14957 3798 14991
rect 4166 14957 4182 14991
rect 3782 14910 4182 14957
rect 3082 14363 3482 14410
rect 3082 14329 3098 14363
rect 3466 14329 3482 14363
rect 3082 14313 3482 14329
rect 3782 14363 4182 14410
rect 3782 14329 3798 14363
rect 4166 14329 4182 14363
rect 3782 14313 4182 14329
rect 3082 14207 3482 14223
rect 3082 14173 3098 14207
rect 3466 14173 3482 14207
rect 3082 14126 3482 14173
rect 3782 14207 4182 14223
rect 3782 14173 3798 14207
rect 4166 14173 4182 14207
rect 3782 14126 4182 14173
rect 3082 13579 3482 13626
rect 3082 13545 3098 13579
rect 3466 13545 3482 13579
rect 3082 13529 3482 13545
rect 3782 13579 4182 13626
rect 3782 13545 3798 13579
rect 4166 13545 4182 13579
rect 3782 13529 4182 13545
rect 3082 13423 3482 13439
rect 3082 13389 3098 13423
rect 3466 13389 3482 13423
rect 3082 13342 3482 13389
rect 3782 13423 4182 13439
rect 3782 13389 3798 13423
rect 4166 13389 4182 13423
rect 3782 13342 4182 13389
rect 3082 12795 3482 12842
rect 3082 12761 3098 12795
rect 3466 12761 3482 12795
rect 3082 12745 3482 12761
rect 3782 12795 4182 12842
rect 3782 12761 3798 12795
rect 4166 12761 4182 12795
rect 3782 12745 4182 12761
rect 3082 12639 3482 12655
rect 3082 12605 3098 12639
rect 3466 12605 3482 12639
rect 3082 12558 3482 12605
rect 3782 12639 4182 12655
rect 3782 12605 3798 12639
rect 4166 12605 4182 12639
rect 3782 12558 4182 12605
rect 3082 12011 3482 12058
rect 3082 11977 3098 12011
rect 3466 11977 3482 12011
rect 3082 11961 3482 11977
rect 3782 12011 4182 12058
rect 3782 11977 3798 12011
rect 4166 11977 4182 12011
rect 3782 11961 4182 11977
rect 3082 11855 3482 11871
rect 3082 11821 3098 11855
rect 3466 11821 3482 11855
rect 3082 11774 3482 11821
rect 3782 11855 4182 11871
rect 3782 11821 3798 11855
rect 4166 11821 4182 11855
rect 3782 11774 4182 11821
rect 3082 11227 3482 11274
rect 3082 11193 3098 11227
rect 3466 11193 3482 11227
rect 3082 11177 3482 11193
rect 3782 11227 4182 11274
rect 3782 11193 3798 11227
rect 4166 11193 4182 11227
rect 3782 11177 4182 11193
rect 3082 11071 3482 11087
rect 3082 11037 3098 11071
rect 3466 11037 3482 11071
rect 3082 10990 3482 11037
rect 3782 11071 4182 11087
rect 3782 11037 3798 11071
rect 4166 11037 4182 11071
rect 3782 10990 4182 11037
rect 3082 10443 3482 10490
rect 3082 10409 3098 10443
rect 3466 10409 3482 10443
rect 3082 10393 3482 10409
rect 3782 10443 4182 10490
rect 3782 10409 3798 10443
rect 4166 10409 4182 10443
rect 3782 10393 4182 10409
rect 3082 10287 3482 10303
rect 3082 10253 3098 10287
rect 3466 10253 3482 10287
rect 3082 10206 3482 10253
rect 3782 10287 4182 10303
rect 3782 10253 3798 10287
rect 4166 10253 4182 10287
rect 3782 10206 4182 10253
rect 3082 9659 3482 9706
rect 3082 9625 3098 9659
rect 3466 9625 3482 9659
rect 3082 9609 3482 9625
rect 3782 9659 4182 9706
rect 3782 9625 3798 9659
rect 4166 9625 4182 9659
rect 3782 9609 4182 9625
rect 3082 9503 3482 9519
rect 3082 9469 3098 9503
rect 3466 9469 3482 9503
rect 3082 9422 3482 9469
rect 3782 9503 4182 9519
rect 3782 9469 3798 9503
rect 4166 9469 4182 9503
rect 3782 9422 4182 9469
rect 3082 8875 3482 8922
rect 3082 8841 3098 8875
rect 3466 8841 3482 8875
rect 3082 8825 3482 8841
rect 3782 8875 4182 8922
rect 3782 8841 3798 8875
rect 4166 8841 4182 8875
rect 3782 8825 4182 8841
rect 3082 8719 3482 8735
rect 3082 8685 3098 8719
rect 3466 8685 3482 8719
rect 3082 8638 3482 8685
rect 3782 8719 4182 8735
rect 3782 8685 3798 8719
rect 4166 8685 4182 8719
rect 3782 8638 4182 8685
rect 3082 8091 3482 8138
rect 3082 8057 3098 8091
rect 3466 8057 3482 8091
rect 3082 8041 3482 8057
rect 3782 8091 4182 8138
rect 3782 8057 3798 8091
rect 4166 8057 4182 8091
rect 3782 8041 4182 8057
rect 3082 7935 3482 7951
rect 3082 7901 3098 7935
rect 3466 7901 3482 7935
rect 3082 7854 3482 7901
rect 3782 7935 4182 7951
rect 3782 7901 3798 7935
rect 4166 7901 4182 7935
rect 3782 7854 4182 7901
rect 3082 7707 3482 7754
rect 3082 7673 3098 7707
rect 3466 7673 3482 7707
rect 3082 7657 3482 7673
rect 3782 7707 4182 7754
rect 3782 7673 3798 7707
rect 4166 7673 4182 7707
rect 3782 7657 4182 7673
rect 5891 19339 6051 19355
rect 5891 19305 5907 19339
rect 6035 19305 6051 19339
rect 5891 19267 6051 19305
rect 6291 19339 6451 19355
rect 6291 19305 6307 19339
rect 6435 19305 6451 19339
rect 6291 19267 6451 19305
rect 6691 19339 6851 19355
rect 6691 19305 6707 19339
rect 6835 19305 6851 19339
rect 6691 19267 6851 19305
rect 7091 19339 7251 19355
rect 7091 19305 7107 19339
rect 7235 19305 7251 19339
rect 7091 19267 7251 19305
rect 7491 19339 7651 19355
rect 7491 19305 7507 19339
rect 7635 19305 7651 19339
rect 7491 19267 7651 19305
rect 7891 19339 8051 19355
rect 7891 19305 7907 19339
rect 8035 19305 8051 19339
rect 7891 19267 8051 19305
rect 8291 19339 8451 19355
rect 8291 19305 8307 19339
rect 8435 19305 8451 19339
rect 8291 19267 8451 19305
rect 8691 19339 8851 19355
rect 8691 19305 8707 19339
rect 8835 19305 8851 19339
rect 8691 19267 8851 19305
rect 9091 19339 9251 19355
rect 9091 19305 9107 19339
rect 9235 19305 9251 19339
rect 9091 19267 9251 19305
rect 9491 19339 9651 19355
rect 9491 19305 9507 19339
rect 9635 19305 9651 19339
rect 9491 19267 9651 19305
rect 9891 19339 10051 19355
rect 9891 19305 9907 19339
rect 10035 19305 10051 19339
rect 9891 19267 10051 19305
rect 10291 19339 10451 19355
rect 10291 19305 10307 19339
rect 10435 19305 10451 19339
rect 10291 19267 10451 19305
rect 10691 19339 10851 19355
rect 10691 19305 10707 19339
rect 10835 19305 10851 19339
rect 10691 19267 10851 19305
rect 11091 19339 11251 19355
rect 11091 19305 11107 19339
rect 11235 19305 11251 19339
rect 11091 19267 11251 19305
rect 11491 19339 11651 19355
rect 11491 19305 11507 19339
rect 11635 19305 11651 19339
rect 11491 19267 11651 19305
rect 11891 19339 12051 19355
rect 11891 19305 11907 19339
rect 12035 19305 12051 19339
rect 11891 19267 12051 19305
rect 5891 18129 6051 18167
rect 5891 18095 5907 18129
rect 6035 18095 6051 18129
rect 5891 18079 6051 18095
rect 6291 18129 6451 18167
rect 6291 18095 6307 18129
rect 6435 18095 6451 18129
rect 6291 18079 6451 18095
rect 6691 18129 6851 18167
rect 6691 18095 6707 18129
rect 6835 18095 6851 18129
rect 6691 18079 6851 18095
rect 7091 18129 7251 18167
rect 7091 18095 7107 18129
rect 7235 18095 7251 18129
rect 7091 18079 7251 18095
rect 7491 18129 7651 18167
rect 7491 18095 7507 18129
rect 7635 18095 7651 18129
rect 7491 18079 7651 18095
rect 7891 18129 8051 18167
rect 7891 18095 7907 18129
rect 8035 18095 8051 18129
rect 7891 18079 8051 18095
rect 8291 18129 8451 18167
rect 8291 18095 8307 18129
rect 8435 18095 8451 18129
rect 8291 18079 8451 18095
rect 8691 18129 8851 18167
rect 8691 18095 8707 18129
rect 8835 18095 8851 18129
rect 8691 18079 8851 18095
rect 9091 18129 9251 18167
rect 9091 18095 9107 18129
rect 9235 18095 9251 18129
rect 9091 18079 9251 18095
rect 9491 18129 9651 18167
rect 9491 18095 9507 18129
rect 9635 18095 9651 18129
rect 9491 18079 9651 18095
rect 9891 18129 10051 18167
rect 9891 18095 9907 18129
rect 10035 18095 10051 18129
rect 9891 18079 10051 18095
rect 10291 18129 10451 18167
rect 10291 18095 10307 18129
rect 10435 18095 10451 18129
rect 10291 18079 10451 18095
rect 10691 18129 10851 18167
rect 10691 18095 10707 18129
rect 10835 18095 10851 18129
rect 10691 18079 10851 18095
rect 11091 18129 11251 18167
rect 11091 18095 11107 18129
rect 11235 18095 11251 18129
rect 11091 18079 11251 18095
rect 11491 18129 11651 18167
rect 11491 18095 11507 18129
rect 11635 18095 11651 18129
rect 11491 18079 11651 18095
rect 11891 18129 12051 18167
rect 11891 18095 11907 18129
rect 12035 18095 12051 18129
rect 11891 18079 12051 18095
rect 5770 17639 5930 17655
rect 5770 17605 5786 17639
rect 5914 17605 5930 17639
rect 5770 17567 5930 17605
rect 6170 17639 6330 17655
rect 6170 17605 6186 17639
rect 6314 17605 6330 17639
rect 6170 17567 6330 17605
rect 6570 17639 6730 17655
rect 6570 17605 6586 17639
rect 6714 17605 6730 17639
rect 6570 17567 6730 17605
rect 6970 17639 7130 17655
rect 6970 17605 6986 17639
rect 7114 17605 7130 17639
rect 6970 17567 7130 17605
rect 7370 17639 7530 17655
rect 7370 17605 7386 17639
rect 7514 17605 7530 17639
rect 7370 17567 7530 17605
rect 7770 17639 7930 17655
rect 7770 17605 7786 17639
rect 7914 17605 7930 17639
rect 7770 17567 7930 17605
rect 8170 17639 8330 17655
rect 8170 17605 8186 17639
rect 8314 17605 8330 17639
rect 8170 17567 8330 17605
rect 8570 17639 8730 17655
rect 8570 17605 8586 17639
rect 8714 17605 8730 17639
rect 8570 17567 8730 17605
rect 9414 17395 9574 17411
rect 9414 17361 9430 17395
rect 9558 17361 9574 17395
rect 9414 17314 9574 17361
rect 9814 17395 9974 17411
rect 9814 17361 9830 17395
rect 9958 17361 9974 17395
rect 9814 17314 9974 17361
rect 9414 17067 9574 17114
rect 9414 17033 9430 17067
rect 9558 17033 9574 17067
rect 9414 17017 9574 17033
rect 9814 17067 9974 17114
rect 9814 17033 9830 17067
rect 9958 17033 9974 17067
rect 9814 17017 9974 17033
rect 10673 17366 10833 17382
rect 10673 17332 10689 17366
rect 10817 17332 10833 17366
rect 10673 17285 10833 17332
rect 11073 17366 11233 17382
rect 11073 17332 11089 17366
rect 11217 17332 11233 17366
rect 11073 17285 11233 17332
rect 11473 17366 11633 17382
rect 11473 17332 11489 17366
rect 11617 17332 11633 17366
rect 11473 17285 11633 17332
rect 11873 17366 12033 17382
rect 11873 17332 11889 17366
rect 12017 17332 12033 17366
rect 11873 17285 12033 17332
rect 10673 17038 10833 17085
rect 10673 17004 10689 17038
rect 10817 17004 10833 17038
rect 10673 16988 10833 17004
rect 11073 17038 11233 17085
rect 11073 17004 11089 17038
rect 11217 17004 11233 17038
rect 11073 16988 11233 17004
rect 11473 17038 11633 17085
rect 11473 17004 11489 17038
rect 11617 17004 11633 17038
rect 11473 16988 11633 17004
rect 11873 17038 12033 17085
rect 11873 17004 11889 17038
rect 12017 17004 12033 17038
rect 11873 16988 12033 17004
rect 5770 16429 5930 16467
rect 5770 16395 5786 16429
rect 5914 16395 5930 16429
rect 5770 16379 5930 16395
rect 6170 16429 6330 16467
rect 6170 16395 6186 16429
rect 6314 16395 6330 16429
rect 6170 16379 6330 16395
rect 6570 16429 6730 16467
rect 6570 16395 6586 16429
rect 6714 16395 6730 16429
rect 6570 16379 6730 16395
rect 6970 16429 7130 16467
rect 6970 16395 6986 16429
rect 7114 16395 7130 16429
rect 6970 16379 7130 16395
rect 7370 16429 7530 16467
rect 7370 16395 7386 16429
rect 7514 16395 7530 16429
rect 7370 16379 7530 16395
rect 7770 16429 7930 16467
rect 7770 16395 7786 16429
rect 7914 16395 7930 16429
rect 7770 16379 7930 16395
rect 8170 16429 8330 16467
rect 8170 16395 8186 16429
rect 8314 16395 8330 16429
rect 8170 16379 8330 16395
rect 8570 16429 8730 16467
rect 8570 16395 8586 16429
rect 8714 16395 8730 16429
rect 8570 16379 8730 16395
rect 5842 15459 5930 15475
rect 5842 15331 5858 15459
rect 5892 15331 5930 15459
rect 5842 15315 5930 15331
rect 7030 15459 7118 15475
rect 7030 15331 7068 15459
rect 7102 15331 7118 15459
rect 7318 15415 7406 15431
rect 7318 15367 7334 15415
rect 7368 15367 7406 15415
rect 7318 15351 7406 15367
rect 8506 15415 8594 15431
rect 8506 15367 8544 15415
rect 8578 15367 8594 15415
rect 8506 15351 8594 15367
rect 7030 15315 7118 15331
rect 7318 15117 7406 15133
rect 5842 15099 5930 15115
rect 5842 14971 5858 15099
rect 5892 14971 5930 15099
rect 5842 14955 5930 14971
rect 7030 15099 7118 15115
rect 7030 14971 7068 15099
rect 7102 14971 7118 15099
rect 7318 15069 7334 15117
rect 7368 15069 7406 15117
rect 7318 15053 7406 15069
rect 8506 15117 8594 15133
rect 8506 15069 8544 15117
rect 8578 15069 8594 15117
rect 8506 15053 8594 15069
rect 7030 14955 7118 14971
rect 7288 14835 7376 14851
rect 5842 14739 5930 14755
rect 5842 14611 5858 14739
rect 5892 14611 5930 14739
rect 5842 14595 5930 14611
rect 7030 14739 7118 14755
rect 7030 14611 7068 14739
rect 7102 14611 7118 14739
rect 7288 14667 7304 14835
rect 7338 14667 7376 14835
rect 7288 14651 7376 14667
rect 8476 14835 8564 14851
rect 8476 14667 8514 14835
rect 8548 14667 8564 14835
rect 8476 14651 8564 14667
rect 7030 14595 7118 14611
rect 7288 14411 7376 14427
rect 5842 14379 5930 14395
rect 5842 14251 5858 14379
rect 5892 14251 5930 14379
rect 5842 14235 5930 14251
rect 7030 14379 7118 14395
rect 7030 14251 7068 14379
rect 7102 14251 7118 14379
rect 7030 14235 7118 14251
rect 7288 14243 7304 14411
rect 7338 14243 7376 14411
rect 7288 14227 7376 14243
rect 8476 14411 8564 14427
rect 8476 14243 8514 14411
rect 8548 14243 8564 14411
rect 8476 14227 8564 14243
rect 8966 15490 9063 15506
rect 8966 15362 8982 15490
rect 9016 15362 9063 15490
rect 8966 15346 9063 15362
rect 9263 15490 9360 15506
rect 9263 15362 9310 15490
rect 9344 15362 9360 15490
rect 9263 15346 9360 15362
rect 8966 15082 9063 15098
rect 8966 14954 8982 15082
rect 9016 14954 9063 15082
rect 8966 14938 9063 14954
rect 9263 15082 9360 15098
rect 9263 14954 9310 15082
rect 9344 14954 9360 15082
rect 9263 14938 9360 14954
rect 8966 14636 9063 14652
rect 8966 14268 8982 14636
rect 9016 14268 9063 14636
rect 8966 14252 9063 14268
rect 9263 14636 9360 14652
rect 9263 14268 9310 14636
rect 9344 14268 9360 14636
rect 9263 14252 9360 14268
rect 9657 15490 9754 15506
rect 9657 15362 9673 15490
rect 9707 15362 9754 15490
rect 9657 15346 9754 15362
rect 9954 15490 10051 15506
rect 9954 15362 10001 15490
rect 10035 15362 10051 15490
rect 9954 15346 10051 15362
rect 9657 15082 9754 15098
rect 9657 14954 9673 15082
rect 9707 14954 9754 15082
rect 9657 14938 9754 14954
rect 9954 15082 10051 15098
rect 9954 14954 10001 15082
rect 10035 14954 10051 15082
rect 9954 14938 10051 14954
rect 9657 14636 9754 14652
rect 9657 14268 9673 14636
rect 9707 14268 9754 14636
rect 9657 14252 9754 14268
rect 9954 14636 10051 14652
rect 9954 14268 10001 14636
rect 10035 14268 10051 14636
rect 9954 14252 10051 14268
rect 11899 15459 11987 15475
rect 10423 15415 10511 15431
rect 10423 15367 10439 15415
rect 10473 15367 10511 15415
rect 10423 15351 10511 15367
rect 11611 15415 11699 15431
rect 11611 15367 11649 15415
rect 11683 15367 11699 15415
rect 11611 15351 11699 15367
rect 11899 15331 11915 15459
rect 11949 15331 11987 15459
rect 11899 15315 11987 15331
rect 13087 15459 13175 15475
rect 13087 15331 13125 15459
rect 13159 15331 13175 15459
rect 13087 15315 13175 15331
rect 10423 15117 10511 15133
rect 10423 15069 10439 15117
rect 10473 15069 10511 15117
rect 10423 15053 10511 15069
rect 11611 15117 11699 15133
rect 11611 15069 11649 15117
rect 11683 15069 11699 15117
rect 11611 15053 11699 15069
rect 11899 15099 11987 15115
rect 11899 14971 11915 15099
rect 11949 14971 11987 15099
rect 11899 14955 11987 14971
rect 13087 15099 13175 15115
rect 13087 14971 13125 15099
rect 13159 14971 13175 15099
rect 13087 14955 13175 14971
rect 10453 14835 10541 14851
rect 10453 14667 10469 14835
rect 10503 14667 10541 14835
rect 10453 14651 10541 14667
rect 11641 14835 11729 14851
rect 11641 14667 11679 14835
rect 11713 14667 11729 14835
rect 11641 14651 11729 14667
rect 11899 14739 11987 14755
rect 11899 14611 11915 14739
rect 11949 14611 11987 14739
rect 11899 14595 11987 14611
rect 13087 14739 13175 14755
rect 13087 14611 13125 14739
rect 13159 14611 13175 14739
rect 13087 14595 13175 14611
rect 10453 14411 10541 14427
rect 10453 14243 10469 14411
rect 10503 14243 10541 14411
rect 10453 14227 10541 14243
rect 11641 14411 11729 14427
rect 11641 14243 11679 14411
rect 11713 14243 11729 14411
rect 11641 14227 11729 14243
rect 11899 14379 11987 14395
rect 11899 14251 11915 14379
rect 11949 14251 11987 14379
rect 11899 14235 11987 14251
rect 13087 14379 13175 14395
rect 13087 14251 13125 14379
rect 13159 14251 13175 14379
rect 13087 14235 13175 14251
rect 5842 13793 5930 13809
rect 5842 13665 5858 13793
rect 5892 13665 5930 13793
rect 5842 13649 5930 13665
rect 7030 13793 7118 13809
rect 7030 13665 7068 13793
rect 7102 13665 7118 13793
rect 7318 13749 7406 13765
rect 7318 13701 7334 13749
rect 7368 13701 7406 13749
rect 7318 13685 7406 13701
rect 8506 13749 8594 13765
rect 8506 13701 8544 13749
rect 8578 13701 8594 13749
rect 8506 13685 8594 13701
rect 7030 13649 7118 13665
rect 7318 13451 7406 13467
rect 5842 13433 5930 13449
rect 5842 13305 5858 13433
rect 5892 13305 5930 13433
rect 5842 13289 5930 13305
rect 7030 13433 7118 13449
rect 7030 13305 7068 13433
rect 7102 13305 7118 13433
rect 7318 13403 7334 13451
rect 7368 13403 7406 13451
rect 7318 13387 7406 13403
rect 8506 13451 8594 13467
rect 8506 13403 8544 13451
rect 8578 13403 8594 13451
rect 8506 13387 8594 13403
rect 7030 13289 7118 13305
rect 7288 13169 7376 13185
rect 5842 13073 5930 13089
rect 5842 12945 5858 13073
rect 5892 12945 5930 13073
rect 5842 12929 5930 12945
rect 7030 13073 7118 13089
rect 7030 12945 7068 13073
rect 7102 12945 7118 13073
rect 7288 13001 7304 13169
rect 7338 13001 7376 13169
rect 7288 12985 7376 13001
rect 8476 13169 8564 13185
rect 8476 13001 8514 13169
rect 8548 13001 8564 13169
rect 8476 12985 8564 13001
rect 7030 12929 7118 12945
rect 7288 12745 7376 12761
rect 5842 12713 5930 12729
rect 5842 12585 5858 12713
rect 5892 12585 5930 12713
rect 5842 12569 5930 12585
rect 7030 12713 7118 12729
rect 7030 12585 7068 12713
rect 7102 12585 7118 12713
rect 7030 12569 7118 12585
rect 7288 12577 7304 12745
rect 7338 12577 7376 12745
rect 7288 12561 7376 12577
rect 8476 12745 8564 12761
rect 8476 12577 8514 12745
rect 8548 12577 8564 12745
rect 8476 12561 8564 12577
rect 8966 13824 9063 13840
rect 8966 13696 8982 13824
rect 9016 13696 9063 13824
rect 8966 13680 9063 13696
rect 9263 13824 9360 13840
rect 9263 13696 9310 13824
rect 9344 13696 9360 13824
rect 9263 13680 9360 13696
rect 8966 13416 9063 13432
rect 8966 13288 8982 13416
rect 9016 13288 9063 13416
rect 8966 13272 9063 13288
rect 9263 13416 9360 13432
rect 9263 13288 9310 13416
rect 9344 13288 9360 13416
rect 9263 13272 9360 13288
rect 8966 12970 9063 12986
rect 8966 12602 8982 12970
rect 9016 12602 9063 12970
rect 8966 12586 9063 12602
rect 9263 12970 9360 12986
rect 9263 12602 9310 12970
rect 9344 12602 9360 12970
rect 9263 12586 9360 12602
rect 9657 13824 9754 13840
rect 9657 13696 9673 13824
rect 9707 13696 9754 13824
rect 9657 13680 9754 13696
rect 9954 13824 10051 13840
rect 9954 13696 10001 13824
rect 10035 13696 10051 13824
rect 9954 13680 10051 13696
rect 9657 13416 9754 13432
rect 9657 13288 9673 13416
rect 9707 13288 9754 13416
rect 9657 13272 9754 13288
rect 9954 13416 10051 13432
rect 9954 13288 10001 13416
rect 10035 13288 10051 13416
rect 9954 13272 10051 13288
rect 9657 12970 9754 12986
rect 9657 12602 9673 12970
rect 9707 12602 9754 12970
rect 9657 12586 9754 12602
rect 9954 12970 10051 12986
rect 9954 12602 10001 12970
rect 10035 12602 10051 12970
rect 9954 12586 10051 12602
rect 11899 13793 11987 13809
rect 10423 13749 10511 13765
rect 10423 13701 10439 13749
rect 10473 13701 10511 13749
rect 10423 13685 10511 13701
rect 11611 13749 11699 13765
rect 11611 13701 11649 13749
rect 11683 13701 11699 13749
rect 11611 13685 11699 13701
rect 11899 13665 11915 13793
rect 11949 13665 11987 13793
rect 11899 13649 11987 13665
rect 13087 13793 13175 13809
rect 13087 13665 13125 13793
rect 13159 13665 13175 13793
rect 13087 13649 13175 13665
rect 10423 13451 10511 13467
rect 10423 13403 10439 13451
rect 10473 13403 10511 13451
rect 10423 13387 10511 13403
rect 11611 13451 11699 13467
rect 11611 13403 11649 13451
rect 11683 13403 11699 13451
rect 11611 13387 11699 13403
rect 11899 13433 11987 13449
rect 11899 13305 11915 13433
rect 11949 13305 11987 13433
rect 11899 13289 11987 13305
rect 13087 13433 13175 13449
rect 13087 13305 13125 13433
rect 13159 13305 13175 13433
rect 13087 13289 13175 13305
rect 10453 13169 10541 13185
rect 10453 13001 10469 13169
rect 10503 13001 10541 13169
rect 10453 12985 10541 13001
rect 11641 13169 11729 13185
rect 11641 13001 11679 13169
rect 11713 13001 11729 13169
rect 11641 12985 11729 13001
rect 11899 13073 11987 13089
rect 11899 12945 11915 13073
rect 11949 12945 11987 13073
rect 11899 12929 11987 12945
rect 13087 13073 13175 13089
rect 13087 12945 13125 13073
rect 13159 12945 13175 13073
rect 13087 12929 13175 12945
rect 10453 12745 10541 12761
rect 10453 12577 10469 12745
rect 10503 12577 10541 12745
rect 10453 12561 10541 12577
rect 11641 12745 11729 12761
rect 11641 12577 11679 12745
rect 11713 12577 11729 12745
rect 11641 12561 11729 12577
rect 11899 12713 11987 12729
rect 11899 12585 11915 12713
rect 11949 12585 11987 12713
rect 11899 12569 11987 12585
rect 13087 12713 13175 12729
rect 13087 12585 13125 12713
rect 13159 12585 13175 12713
rect 13087 12569 13175 12585
rect 5842 12127 5930 12143
rect 5842 11999 5858 12127
rect 5892 11999 5930 12127
rect 5842 11983 5930 11999
rect 7030 12127 7118 12143
rect 7030 11999 7068 12127
rect 7102 11999 7118 12127
rect 7318 12083 7406 12099
rect 7318 12035 7334 12083
rect 7368 12035 7406 12083
rect 7318 12019 7406 12035
rect 8506 12083 8594 12099
rect 8506 12035 8544 12083
rect 8578 12035 8594 12083
rect 8506 12019 8594 12035
rect 7030 11983 7118 11999
rect 7318 11785 7406 11801
rect 5842 11767 5930 11783
rect 5842 11639 5858 11767
rect 5892 11639 5930 11767
rect 5842 11623 5930 11639
rect 7030 11767 7118 11783
rect 7030 11639 7068 11767
rect 7102 11639 7118 11767
rect 7318 11737 7334 11785
rect 7368 11737 7406 11785
rect 7318 11721 7406 11737
rect 8506 11785 8594 11801
rect 8506 11737 8544 11785
rect 8578 11737 8594 11785
rect 8506 11721 8594 11737
rect 7030 11623 7118 11639
rect 7288 11503 7376 11519
rect 5842 11407 5930 11423
rect 5842 11279 5858 11407
rect 5892 11279 5930 11407
rect 5842 11263 5930 11279
rect 7030 11407 7118 11423
rect 7030 11279 7068 11407
rect 7102 11279 7118 11407
rect 7288 11335 7304 11503
rect 7338 11335 7376 11503
rect 7288 11319 7376 11335
rect 8476 11503 8564 11519
rect 8476 11335 8514 11503
rect 8548 11335 8564 11503
rect 8476 11319 8564 11335
rect 7030 11263 7118 11279
rect 7288 11079 7376 11095
rect 5842 11047 5930 11063
rect 5842 10919 5858 11047
rect 5892 10919 5930 11047
rect 5842 10903 5930 10919
rect 7030 11047 7118 11063
rect 7030 10919 7068 11047
rect 7102 10919 7118 11047
rect 7030 10903 7118 10919
rect 7288 10911 7304 11079
rect 7338 10911 7376 11079
rect 7288 10895 7376 10911
rect 8476 11079 8564 11095
rect 8476 10911 8514 11079
rect 8548 10911 8564 11079
rect 8476 10895 8564 10911
rect 8966 12158 9063 12174
rect 8966 12030 8982 12158
rect 9016 12030 9063 12158
rect 8966 12014 9063 12030
rect 9263 12158 9360 12174
rect 9263 12030 9310 12158
rect 9344 12030 9360 12158
rect 9263 12014 9360 12030
rect 8966 11750 9063 11766
rect 8966 11622 8982 11750
rect 9016 11622 9063 11750
rect 8966 11606 9063 11622
rect 9263 11750 9360 11766
rect 9263 11622 9310 11750
rect 9344 11622 9360 11750
rect 9263 11606 9360 11622
rect 8966 11304 9063 11320
rect 8966 10936 8982 11304
rect 9016 10936 9063 11304
rect 8966 10920 9063 10936
rect 9263 11304 9360 11320
rect 9263 10936 9310 11304
rect 9344 10936 9360 11304
rect 9263 10920 9360 10936
rect 9657 12158 9754 12174
rect 9657 12030 9673 12158
rect 9707 12030 9754 12158
rect 9657 12014 9754 12030
rect 9954 12158 10051 12174
rect 9954 12030 10001 12158
rect 10035 12030 10051 12158
rect 9954 12014 10051 12030
rect 9657 11750 9754 11766
rect 9657 11622 9673 11750
rect 9707 11622 9754 11750
rect 9657 11606 9754 11622
rect 9954 11750 10051 11766
rect 9954 11622 10001 11750
rect 10035 11622 10051 11750
rect 9954 11606 10051 11622
rect 9657 11304 9754 11320
rect 9657 10936 9673 11304
rect 9707 10936 9754 11304
rect 9657 10920 9754 10936
rect 9954 11304 10051 11320
rect 9954 10936 10001 11304
rect 10035 10936 10051 11304
rect 9954 10920 10051 10936
rect 11899 12127 11987 12143
rect 10423 12083 10511 12099
rect 10423 12035 10439 12083
rect 10473 12035 10511 12083
rect 10423 12019 10511 12035
rect 11611 12083 11699 12099
rect 11611 12035 11649 12083
rect 11683 12035 11699 12083
rect 11611 12019 11699 12035
rect 11899 11999 11915 12127
rect 11949 11999 11987 12127
rect 11899 11983 11987 11999
rect 13087 12127 13175 12143
rect 13087 11999 13125 12127
rect 13159 11999 13175 12127
rect 13087 11983 13175 11999
rect 10423 11785 10511 11801
rect 10423 11737 10439 11785
rect 10473 11737 10511 11785
rect 10423 11721 10511 11737
rect 11611 11785 11699 11801
rect 11611 11737 11649 11785
rect 11683 11737 11699 11785
rect 11611 11721 11699 11737
rect 11899 11767 11987 11783
rect 11899 11639 11915 11767
rect 11949 11639 11987 11767
rect 11899 11623 11987 11639
rect 13087 11767 13175 11783
rect 13087 11639 13125 11767
rect 13159 11639 13175 11767
rect 13087 11623 13175 11639
rect 10453 11503 10541 11519
rect 10453 11335 10469 11503
rect 10503 11335 10541 11503
rect 10453 11319 10541 11335
rect 11641 11503 11729 11519
rect 11641 11335 11679 11503
rect 11713 11335 11729 11503
rect 11641 11319 11729 11335
rect 11899 11407 11987 11423
rect 11899 11279 11915 11407
rect 11949 11279 11987 11407
rect 11899 11263 11987 11279
rect 13087 11407 13175 11423
rect 13087 11279 13125 11407
rect 13159 11279 13175 11407
rect 13087 11263 13175 11279
rect 10453 11079 10541 11095
rect 10453 10911 10469 11079
rect 10503 10911 10541 11079
rect 10453 10895 10541 10911
rect 11641 11079 11729 11095
rect 11641 10911 11679 11079
rect 11713 10911 11729 11079
rect 11641 10895 11729 10911
rect 11899 11047 11987 11063
rect 11899 10919 11915 11047
rect 11949 10919 11987 11047
rect 11899 10903 11987 10919
rect 13087 11047 13175 11063
rect 13087 10919 13125 11047
rect 13159 10919 13175 11047
rect 13087 10903 13175 10919
rect 5842 10461 5930 10477
rect 5842 10333 5858 10461
rect 5892 10333 5930 10461
rect 5842 10317 5930 10333
rect 7030 10461 7118 10477
rect 7030 10333 7068 10461
rect 7102 10333 7118 10461
rect 7318 10417 7406 10433
rect 7318 10369 7334 10417
rect 7368 10369 7406 10417
rect 7318 10353 7406 10369
rect 8506 10417 8594 10433
rect 8506 10369 8544 10417
rect 8578 10369 8594 10417
rect 8506 10353 8594 10369
rect 7030 10317 7118 10333
rect 7318 10119 7406 10135
rect 5842 10101 5930 10117
rect 5842 9973 5858 10101
rect 5892 9973 5930 10101
rect 5842 9957 5930 9973
rect 7030 10101 7118 10117
rect 7030 9973 7068 10101
rect 7102 9973 7118 10101
rect 7318 10071 7334 10119
rect 7368 10071 7406 10119
rect 7318 10055 7406 10071
rect 8506 10119 8594 10135
rect 8506 10071 8544 10119
rect 8578 10071 8594 10119
rect 8506 10055 8594 10071
rect 7030 9957 7118 9973
rect 7288 9837 7376 9853
rect 5842 9741 5930 9757
rect 5842 9613 5858 9741
rect 5892 9613 5930 9741
rect 5842 9597 5930 9613
rect 7030 9741 7118 9757
rect 7030 9613 7068 9741
rect 7102 9613 7118 9741
rect 7288 9669 7304 9837
rect 7338 9669 7376 9837
rect 7288 9653 7376 9669
rect 8476 9837 8564 9853
rect 8476 9669 8514 9837
rect 8548 9669 8564 9837
rect 8476 9653 8564 9669
rect 7030 9597 7118 9613
rect 7288 9413 7376 9429
rect 5842 9381 5930 9397
rect 5842 9253 5858 9381
rect 5892 9253 5930 9381
rect 5842 9237 5930 9253
rect 7030 9381 7118 9397
rect 7030 9253 7068 9381
rect 7102 9253 7118 9381
rect 7030 9237 7118 9253
rect 7288 9245 7304 9413
rect 7338 9245 7376 9413
rect 7288 9229 7376 9245
rect 8476 9413 8564 9429
rect 8476 9245 8514 9413
rect 8548 9245 8564 9413
rect 8476 9229 8564 9245
rect 8966 10492 9063 10508
rect 8966 10364 8982 10492
rect 9016 10364 9063 10492
rect 8966 10348 9063 10364
rect 9263 10492 9360 10508
rect 9263 10364 9310 10492
rect 9344 10364 9360 10492
rect 9263 10348 9360 10364
rect 8966 10084 9063 10100
rect 8966 9956 8982 10084
rect 9016 9956 9063 10084
rect 8966 9940 9063 9956
rect 9263 10084 9360 10100
rect 9263 9956 9310 10084
rect 9344 9956 9360 10084
rect 9263 9940 9360 9956
rect 8966 9638 9063 9654
rect 8966 9270 8982 9638
rect 9016 9270 9063 9638
rect 8966 9254 9063 9270
rect 9263 9638 9360 9654
rect 9263 9270 9310 9638
rect 9344 9270 9360 9638
rect 9263 9254 9360 9270
rect 9657 10492 9754 10508
rect 9657 10364 9673 10492
rect 9707 10364 9754 10492
rect 9657 10348 9754 10364
rect 9954 10492 10051 10508
rect 9954 10364 10001 10492
rect 10035 10364 10051 10492
rect 9954 10348 10051 10364
rect 9657 10084 9754 10100
rect 9657 9956 9673 10084
rect 9707 9956 9754 10084
rect 9657 9940 9754 9956
rect 9954 10084 10051 10100
rect 9954 9956 10001 10084
rect 10035 9956 10051 10084
rect 9954 9940 10051 9956
rect 9657 9638 9754 9654
rect 9657 9270 9673 9638
rect 9707 9270 9754 9638
rect 9657 9254 9754 9270
rect 9954 9638 10051 9654
rect 9954 9270 10001 9638
rect 10035 9270 10051 9638
rect 9954 9254 10051 9270
rect 11899 10461 11987 10477
rect 10423 10417 10511 10433
rect 10423 10369 10439 10417
rect 10473 10369 10511 10417
rect 10423 10353 10511 10369
rect 11611 10417 11699 10433
rect 11611 10369 11649 10417
rect 11683 10369 11699 10417
rect 11611 10353 11699 10369
rect 11899 10333 11915 10461
rect 11949 10333 11987 10461
rect 11899 10317 11987 10333
rect 13087 10461 13175 10477
rect 13087 10333 13125 10461
rect 13159 10333 13175 10461
rect 13087 10317 13175 10333
rect 10423 10119 10511 10135
rect 10423 10071 10439 10119
rect 10473 10071 10511 10119
rect 10423 10055 10511 10071
rect 11611 10119 11699 10135
rect 11611 10071 11649 10119
rect 11683 10071 11699 10119
rect 11611 10055 11699 10071
rect 11899 10101 11987 10117
rect 11899 9973 11915 10101
rect 11949 9973 11987 10101
rect 11899 9957 11987 9973
rect 13087 10101 13175 10117
rect 13087 9973 13125 10101
rect 13159 9973 13175 10101
rect 13087 9957 13175 9973
rect 10453 9837 10541 9853
rect 10453 9669 10469 9837
rect 10503 9669 10541 9837
rect 10453 9653 10541 9669
rect 11641 9837 11729 9853
rect 11641 9669 11679 9837
rect 11713 9669 11729 9837
rect 11641 9653 11729 9669
rect 11899 9741 11987 9757
rect 11899 9613 11915 9741
rect 11949 9613 11987 9741
rect 11899 9597 11987 9613
rect 13087 9741 13175 9757
rect 13087 9613 13125 9741
rect 13159 9613 13175 9741
rect 13087 9597 13175 9613
rect 10453 9413 10541 9429
rect 10453 9245 10469 9413
rect 10503 9245 10541 9413
rect 10453 9229 10541 9245
rect 11641 9413 11729 9429
rect 11641 9245 11679 9413
rect 11713 9245 11729 9413
rect 11641 9229 11729 9245
rect 11899 9381 11987 9397
rect 11899 9253 11915 9381
rect 11949 9253 11987 9381
rect 11899 9237 11987 9253
rect 13087 9381 13175 9397
rect 13087 9253 13125 9381
rect 13159 9253 13175 9381
rect 13087 9237 13175 9253
rect 5842 8795 5930 8811
rect 5842 8667 5858 8795
rect 5892 8667 5930 8795
rect 5842 8651 5930 8667
rect 7030 8795 7118 8811
rect 7030 8667 7068 8795
rect 7102 8667 7118 8795
rect 7318 8751 7406 8767
rect 7318 8703 7334 8751
rect 7368 8703 7406 8751
rect 7318 8687 7406 8703
rect 8506 8751 8594 8767
rect 8506 8703 8544 8751
rect 8578 8703 8594 8751
rect 8506 8687 8594 8703
rect 7030 8651 7118 8667
rect 7318 8453 7406 8469
rect 5842 8435 5930 8451
rect 5842 8307 5858 8435
rect 5892 8307 5930 8435
rect 5842 8291 5930 8307
rect 7030 8435 7118 8451
rect 7030 8307 7068 8435
rect 7102 8307 7118 8435
rect 7318 8405 7334 8453
rect 7368 8405 7406 8453
rect 7318 8389 7406 8405
rect 8506 8453 8594 8469
rect 8506 8405 8544 8453
rect 8578 8405 8594 8453
rect 8506 8389 8594 8405
rect 7030 8291 7118 8307
rect 7288 8171 7376 8187
rect 5842 8075 5930 8091
rect 5842 7947 5858 8075
rect 5892 7947 5930 8075
rect 5842 7931 5930 7947
rect 7030 8075 7118 8091
rect 7030 7947 7068 8075
rect 7102 7947 7118 8075
rect 7288 8003 7304 8171
rect 7338 8003 7376 8171
rect 7288 7987 7376 8003
rect 8476 8171 8564 8187
rect 8476 8003 8514 8171
rect 8548 8003 8564 8171
rect 8476 7987 8564 8003
rect 7030 7931 7118 7947
rect 7288 7747 7376 7763
rect 5842 7715 5930 7731
rect 5842 7587 5858 7715
rect 5892 7587 5930 7715
rect 5842 7571 5930 7587
rect 7030 7715 7118 7731
rect 7030 7587 7068 7715
rect 7102 7587 7118 7715
rect 7030 7571 7118 7587
rect 7288 7579 7304 7747
rect 7338 7579 7376 7747
rect 7288 7563 7376 7579
rect 8476 7747 8564 7763
rect 8476 7579 8514 7747
rect 8548 7579 8564 7747
rect 8476 7563 8564 7579
rect 8966 8826 9063 8842
rect 8966 8698 8982 8826
rect 9016 8698 9063 8826
rect 8966 8682 9063 8698
rect 9263 8826 9360 8842
rect 9263 8698 9310 8826
rect 9344 8698 9360 8826
rect 9263 8682 9360 8698
rect 8966 8418 9063 8434
rect 8966 8290 8982 8418
rect 9016 8290 9063 8418
rect 8966 8274 9063 8290
rect 9263 8418 9360 8434
rect 9263 8290 9310 8418
rect 9344 8290 9360 8418
rect 9263 8274 9360 8290
rect 8966 7972 9063 7988
rect 8966 7604 8982 7972
rect 9016 7604 9063 7972
rect 8966 7588 9063 7604
rect 9263 7972 9360 7988
rect 9263 7604 9310 7972
rect 9344 7604 9360 7972
rect 9263 7588 9360 7604
rect 9657 8826 9754 8842
rect 9657 8698 9673 8826
rect 9707 8698 9754 8826
rect 9657 8682 9754 8698
rect 9954 8826 10051 8842
rect 9954 8698 10001 8826
rect 10035 8698 10051 8826
rect 9954 8682 10051 8698
rect 9657 8418 9754 8434
rect 9657 8290 9673 8418
rect 9707 8290 9754 8418
rect 9657 8274 9754 8290
rect 9954 8418 10051 8434
rect 9954 8290 10001 8418
rect 10035 8290 10051 8418
rect 9954 8274 10051 8290
rect 9657 7972 9754 7988
rect 9657 7604 9673 7972
rect 9707 7604 9754 7972
rect 9657 7588 9754 7604
rect 9954 7972 10051 7988
rect 9954 7604 10001 7972
rect 10035 7604 10051 7972
rect 9954 7588 10051 7604
rect 11899 8795 11987 8811
rect 10423 8751 10511 8767
rect 10423 8703 10439 8751
rect 10473 8703 10511 8751
rect 10423 8687 10511 8703
rect 11611 8751 11699 8767
rect 11611 8703 11649 8751
rect 11683 8703 11699 8751
rect 11611 8687 11699 8703
rect 11899 8667 11915 8795
rect 11949 8667 11987 8795
rect 11899 8651 11987 8667
rect 13087 8795 13175 8811
rect 13087 8667 13125 8795
rect 13159 8667 13175 8795
rect 13087 8651 13175 8667
rect 10423 8453 10511 8469
rect 10423 8405 10439 8453
rect 10473 8405 10511 8453
rect 10423 8389 10511 8405
rect 11611 8453 11699 8469
rect 11611 8405 11649 8453
rect 11683 8405 11699 8453
rect 11611 8389 11699 8405
rect 11899 8435 11987 8451
rect 11899 8307 11915 8435
rect 11949 8307 11987 8435
rect 11899 8291 11987 8307
rect 13087 8435 13175 8451
rect 13087 8307 13125 8435
rect 13159 8307 13175 8435
rect 13087 8291 13175 8307
rect 10453 8171 10541 8187
rect 10453 8003 10469 8171
rect 10503 8003 10541 8171
rect 10453 7987 10541 8003
rect 11641 8171 11729 8187
rect 11641 8003 11679 8171
rect 11713 8003 11729 8171
rect 11641 7987 11729 8003
rect 11899 8075 11987 8091
rect 11899 7947 11915 8075
rect 11949 7947 11987 8075
rect 11899 7931 11987 7947
rect 13087 8075 13175 8091
rect 13087 7947 13125 8075
rect 13159 7947 13175 8075
rect 13087 7931 13175 7947
rect 10453 7747 10541 7763
rect 10453 7579 10469 7747
rect 10503 7579 10541 7747
rect 10453 7563 10541 7579
rect 11641 7747 11729 7763
rect 11641 7579 11679 7747
rect 11713 7579 11729 7747
rect 11641 7563 11729 7579
rect 11899 7715 11987 7731
rect 11899 7587 11915 7715
rect 11949 7587 11987 7715
rect 11899 7571 11987 7587
rect 13087 7715 13175 7731
rect 13087 7587 13125 7715
rect 13159 7587 13175 7715
rect 13087 7571 13175 7587
rect 15101 17766 15171 17782
rect 15101 17732 15117 17766
rect 15155 17732 15171 17766
rect 15101 17685 15171 17732
rect 15101 15918 15171 15965
rect 15101 15884 15117 15918
rect 15155 15884 15171 15918
rect 15101 15868 15171 15884
rect 16150 17434 16238 17450
rect 16150 17288 16166 17434
rect 16200 17288 16238 17434
rect 16150 17272 16238 17288
rect 17438 17434 17526 17450
rect 17438 17288 17476 17434
rect 17510 17288 17526 17434
rect 17438 17272 17526 17288
rect 16150 17064 16238 17080
rect 16150 16918 16166 17064
rect 16200 16918 16238 17064
rect 16150 16902 16238 16918
rect 17438 17064 17526 17080
rect 17438 16918 17476 17064
rect 17510 16918 17526 17064
rect 17438 16902 17526 16918
rect 16532 16728 17152 16744
rect 16532 16694 16548 16728
rect 17136 16694 17152 16728
rect 16532 16656 17152 16694
rect 17420 16656 17630 16672
rect 17420 16622 17436 16656
rect 17614 16622 17630 16656
rect 17420 16584 17630 16622
rect 17420 16382 17630 16420
rect 17420 16348 17436 16382
rect 17614 16348 17630 16382
rect 17420 16332 17630 16348
rect 16532 16274 17152 16312
rect 16532 16240 16548 16274
rect 17136 16240 17152 16274
rect 16532 16224 17152 16240
rect 14885 13440 14982 13456
rect 14885 12694 14901 13440
rect 14935 12694 14982 13440
rect 14885 12678 14982 12694
rect 15160 13440 15257 13456
rect 15160 12694 15207 13440
rect 15241 12694 15257 13440
rect 15160 12678 15257 12694
rect 15385 13440 15482 13456
rect 15385 12694 15401 13440
rect 15435 12694 15482 13440
rect 15385 12678 15482 12694
rect 15660 13440 15757 13456
rect 15660 12694 15707 13440
rect 15741 12694 15757 13440
rect 15660 12678 15757 12694
rect 15885 13440 15982 13456
rect 15885 12694 15901 13440
rect 15935 12694 15982 13440
rect 15885 12678 15982 12694
rect 16160 13440 16257 13456
rect 16160 12694 16207 13440
rect 16241 12694 16257 13440
rect 16160 12678 16257 12694
rect 16385 13440 16482 13456
rect 16385 12694 16401 13440
rect 16435 12694 16482 13440
rect 16385 12678 16482 12694
rect 16660 13440 16757 13456
rect 16660 12694 16707 13440
rect 16741 12694 16757 13440
rect 16660 12678 16757 12694
rect 16885 13440 16982 13456
rect 16885 12694 16901 13440
rect 16935 12694 16982 13440
rect 16885 12678 16982 12694
rect 17160 13440 17257 13456
rect 17160 12694 17207 13440
rect 17241 12694 17257 13440
rect 17160 12678 17257 12694
rect 17385 13440 17482 13456
rect 17385 12694 17401 13440
rect 17435 12694 17482 13440
rect 17385 12678 17482 12694
rect 17660 13440 17757 13456
rect 17660 12694 17707 13440
rect 17741 12694 17757 13440
rect 17660 12678 17757 12694
rect 14548 11746 14834 11762
rect 14548 11712 14564 11746
rect 14818 11712 14834 11746
rect 14548 11674 14834 11712
rect 14548 10598 14834 10636
rect 14548 10564 14564 10598
rect 14818 10564 14834 10598
rect 14548 10548 14834 10564
rect 14548 10490 14834 10506
rect 14548 10456 14564 10490
rect 14818 10456 14834 10490
rect 14548 10418 14834 10456
rect 14548 9342 14834 9380
rect 14548 9308 14564 9342
rect 14818 9308 14834 9342
rect 14548 9292 14834 9308
rect 16989 11285 17086 11301
rect 16989 11243 17005 11285
rect 17039 11243 17086 11285
rect 16989 11227 17086 11243
rect 18120 11285 18217 11301
rect 18120 11243 18167 11285
rect 18201 11243 18217 11285
rect 18120 11227 18217 11243
rect 16932 10218 17029 10234
rect 16932 9996 16948 10218
rect 16982 9996 17029 10218
rect 16932 9980 17029 9996
rect 18243 10218 18340 10234
rect 18243 9996 18290 10218
rect 18324 9996 18340 10218
rect 18243 9980 18340 9996
rect 16932 9618 17029 9634
rect 16932 9396 16948 9618
rect 16982 9396 17029 9618
rect 16932 9380 17029 9396
rect 18243 9618 18340 9634
rect 18243 9396 18290 9618
rect 18324 9396 18340 9618
rect 18243 9380 18340 9396
rect 14522 8670 14654 8686
rect 14522 8636 14538 8670
rect 14638 8636 14654 8670
rect 14522 8598 14654 8636
rect 14922 8670 15054 8686
rect 14922 8636 14938 8670
rect 15038 8636 15054 8670
rect 14922 8598 15054 8636
rect 15322 8670 15454 8686
rect 15322 8636 15338 8670
rect 15438 8636 15454 8670
rect 15322 8598 15454 8636
rect 15722 8670 15854 8686
rect 15722 8636 15738 8670
rect 15838 8636 15854 8670
rect 15722 8598 15854 8636
rect 16122 8670 16254 8686
rect 16122 8636 16138 8670
rect 16238 8636 16254 8670
rect 16122 8598 16254 8636
rect 16522 8670 16654 8686
rect 16522 8636 16538 8670
rect 16638 8636 16654 8670
rect 16522 8598 16654 8636
rect 16922 8670 17054 8686
rect 16922 8636 16938 8670
rect 17038 8636 17054 8670
rect 16922 8598 17054 8636
rect 17322 8670 17454 8686
rect 17322 8636 17338 8670
rect 17438 8636 17454 8670
rect 17322 8598 17454 8636
rect 17722 8670 17854 8686
rect 17722 8636 17738 8670
rect 17838 8636 17854 8670
rect 17722 8598 17854 8636
rect 18122 8670 18254 8686
rect 18122 8636 18138 8670
rect 18238 8636 18254 8670
rect 18122 8598 18254 8636
rect 14522 7540 14654 7578
rect 14522 7506 14538 7540
rect 14638 7506 14654 7540
rect 14522 7490 14654 7506
rect 14922 7540 15054 7578
rect 14922 7506 14938 7540
rect 15038 7506 15054 7540
rect 14922 7490 15054 7506
rect 15322 7540 15454 7578
rect 15322 7506 15338 7540
rect 15438 7506 15454 7540
rect 15322 7490 15454 7506
rect 15722 7540 15854 7578
rect 15722 7506 15738 7540
rect 15838 7506 15854 7540
rect 15722 7490 15854 7506
rect 16122 7540 16254 7578
rect 16122 7506 16138 7540
rect 16238 7506 16254 7540
rect 16122 7490 16254 7506
rect 16522 7540 16654 7578
rect 16522 7506 16538 7540
rect 16638 7506 16654 7540
rect 16522 7490 16654 7506
rect 16922 7540 17054 7578
rect 16922 7506 16938 7540
rect 17038 7506 17054 7540
rect 16922 7490 17054 7506
rect 17322 7540 17454 7578
rect 17322 7506 17338 7540
rect 17438 7506 17454 7540
rect 17322 7490 17454 7506
rect 17722 7540 17854 7578
rect 17722 7506 17738 7540
rect 17838 7506 17854 7540
rect 17722 7490 17854 7506
rect 18122 7540 18254 7578
rect 18122 7506 18138 7540
rect 18238 7506 18254 7540
rect 18122 7490 18254 7506
<< polycont >>
rect -153 18799 -119 18967
rect 457 18799 491 18967
rect -153 18383 -119 18551
rect 457 18383 491 18551
rect -153 17967 -119 18135
rect 457 17967 491 18135
rect -153 17551 -119 17719
rect 457 17551 491 17719
rect -153 17135 -119 17303
rect 457 17135 491 17303
rect -153 16719 -119 16887
rect 457 16719 491 16887
rect -153 16303 -119 16471
rect 457 16303 491 16471
rect -153 15887 -119 16055
rect 457 15887 491 16055
rect 1402 19245 1770 19279
rect 2102 19245 2470 19279
rect 1402 19017 1770 19051
rect 2102 19017 2470 19051
rect 1402 18861 1770 18895
rect 2102 18861 2470 18895
rect 1402 18233 1770 18267
rect 2102 18233 2470 18267
rect 1402 18077 1770 18111
rect 2102 18077 2470 18111
rect 1402 17449 1770 17483
rect 2102 17449 2470 17483
rect 1402 17293 1770 17327
rect 2102 17293 2470 17327
rect 1402 16665 1770 16699
rect 2102 16665 2470 16699
rect 1402 16509 1770 16543
rect 2102 16509 2470 16543
rect 1402 15881 1770 15915
rect 2102 15881 2470 15915
rect 1402 15725 1770 15759
rect 2102 15725 2470 15759
rect 1402 15497 1770 15531
rect 2102 15497 2470 15531
rect 70 14651 238 14685
rect 486 14651 654 14685
rect 902 14651 1070 14685
rect 1318 14651 1486 14685
rect 1734 14651 1902 14685
rect 2150 14651 2318 14685
rect 70 14041 238 14075
rect 486 14041 654 14075
rect 902 14041 1070 14075
rect 1318 14041 1486 14075
rect 1734 14041 1902 14075
rect 2150 14041 2318 14075
rect 675 13767 1643 13801
rect 675 13457 1643 13491
rect -244 12596 -210 12664
rect 284 12596 318 12664
rect 392 12596 426 12664
rect 920 12596 954 12664
rect 1028 12596 1062 12664
rect 1556 12596 1590 12664
rect 1664 12596 1698 12664
rect 2192 12596 2226 12664
rect 795 11946 2157 11980
rect 795 11642 2157 11676
rect 417 11044 939 11078
rect 1411 11038 2179 11072
rect 1411 10810 2179 10844
rect 1337 10646 2181 10680
rect 417 10230 939 10264
rect 1337 10044 2181 10078
rect 1171 9299 1539 9333
rect 1871 9299 2239 9333
rect 1171 8671 1539 8705
rect 1871 8671 2239 8705
rect 1171 8515 1539 8549
rect 1871 8515 2239 8549
rect 1171 7887 1539 7921
rect 1871 7887 2239 7921
rect 3098 19261 3466 19295
rect 3798 19261 4166 19295
rect 3098 19033 3466 19067
rect 3798 19033 4166 19067
rect 3098 18877 3466 18911
rect 3798 18877 4166 18911
rect 3098 18249 3466 18283
rect 3798 18249 4166 18283
rect 3098 18093 3466 18127
rect 3798 18093 4166 18127
rect 3098 17465 3466 17499
rect 3798 17465 4166 17499
rect 3098 17309 3466 17343
rect 3798 17309 4166 17343
rect 3098 16681 3466 16715
rect 3798 16681 4166 16715
rect 3098 16525 3466 16559
rect 3798 16525 4166 16559
rect 3098 15897 3466 15931
rect 3798 15897 4166 15931
rect 3098 15741 3466 15775
rect 3798 15741 4166 15775
rect 3098 15113 3466 15147
rect 3798 15113 4166 15147
rect 3098 14957 3466 14991
rect 3798 14957 4166 14991
rect 3098 14329 3466 14363
rect 3798 14329 4166 14363
rect 3098 14173 3466 14207
rect 3798 14173 4166 14207
rect 3098 13545 3466 13579
rect 3798 13545 4166 13579
rect 3098 13389 3466 13423
rect 3798 13389 4166 13423
rect 3098 12761 3466 12795
rect 3798 12761 4166 12795
rect 3098 12605 3466 12639
rect 3798 12605 4166 12639
rect 3098 11977 3466 12011
rect 3798 11977 4166 12011
rect 3098 11821 3466 11855
rect 3798 11821 4166 11855
rect 3098 11193 3466 11227
rect 3798 11193 4166 11227
rect 3098 11037 3466 11071
rect 3798 11037 4166 11071
rect 3098 10409 3466 10443
rect 3798 10409 4166 10443
rect 3098 10253 3466 10287
rect 3798 10253 4166 10287
rect 3098 9625 3466 9659
rect 3798 9625 4166 9659
rect 3098 9469 3466 9503
rect 3798 9469 4166 9503
rect 3098 8841 3466 8875
rect 3798 8841 4166 8875
rect 3098 8685 3466 8719
rect 3798 8685 4166 8719
rect 3098 8057 3466 8091
rect 3798 8057 4166 8091
rect 3098 7901 3466 7935
rect 3798 7901 4166 7935
rect 3098 7673 3466 7707
rect 3798 7673 4166 7707
rect 5907 19305 6035 19339
rect 6307 19305 6435 19339
rect 6707 19305 6835 19339
rect 7107 19305 7235 19339
rect 7507 19305 7635 19339
rect 7907 19305 8035 19339
rect 8307 19305 8435 19339
rect 8707 19305 8835 19339
rect 9107 19305 9235 19339
rect 9507 19305 9635 19339
rect 9907 19305 10035 19339
rect 10307 19305 10435 19339
rect 10707 19305 10835 19339
rect 11107 19305 11235 19339
rect 11507 19305 11635 19339
rect 11907 19305 12035 19339
rect 5907 18095 6035 18129
rect 6307 18095 6435 18129
rect 6707 18095 6835 18129
rect 7107 18095 7235 18129
rect 7507 18095 7635 18129
rect 7907 18095 8035 18129
rect 8307 18095 8435 18129
rect 8707 18095 8835 18129
rect 9107 18095 9235 18129
rect 9507 18095 9635 18129
rect 9907 18095 10035 18129
rect 10307 18095 10435 18129
rect 10707 18095 10835 18129
rect 11107 18095 11235 18129
rect 11507 18095 11635 18129
rect 11907 18095 12035 18129
rect 5786 17605 5914 17639
rect 6186 17605 6314 17639
rect 6586 17605 6714 17639
rect 6986 17605 7114 17639
rect 7386 17605 7514 17639
rect 7786 17605 7914 17639
rect 8186 17605 8314 17639
rect 8586 17605 8714 17639
rect 9430 17361 9558 17395
rect 9830 17361 9958 17395
rect 9430 17033 9558 17067
rect 9830 17033 9958 17067
rect 10689 17332 10817 17366
rect 11089 17332 11217 17366
rect 11489 17332 11617 17366
rect 11889 17332 12017 17366
rect 10689 17004 10817 17038
rect 11089 17004 11217 17038
rect 11489 17004 11617 17038
rect 11889 17004 12017 17038
rect 5786 16395 5914 16429
rect 6186 16395 6314 16429
rect 6586 16395 6714 16429
rect 6986 16395 7114 16429
rect 7386 16395 7514 16429
rect 7786 16395 7914 16429
rect 8186 16395 8314 16429
rect 8586 16395 8714 16429
rect 5858 15331 5892 15459
rect 7068 15331 7102 15459
rect 7334 15367 7368 15415
rect 8544 15367 8578 15415
rect 5858 14971 5892 15099
rect 7068 14971 7102 15099
rect 7334 15069 7368 15117
rect 8544 15069 8578 15117
rect 5858 14611 5892 14739
rect 7068 14611 7102 14739
rect 7304 14667 7338 14835
rect 8514 14667 8548 14835
rect 5858 14251 5892 14379
rect 7068 14251 7102 14379
rect 7304 14243 7338 14411
rect 8514 14243 8548 14411
rect 8982 15362 9016 15490
rect 9310 15362 9344 15490
rect 8982 14954 9016 15082
rect 9310 14954 9344 15082
rect 8982 14268 9016 14636
rect 9310 14268 9344 14636
rect 9673 15362 9707 15490
rect 10001 15362 10035 15490
rect 9673 14954 9707 15082
rect 10001 14954 10035 15082
rect 9673 14268 9707 14636
rect 10001 14268 10035 14636
rect 10439 15367 10473 15415
rect 11649 15367 11683 15415
rect 11915 15331 11949 15459
rect 13125 15331 13159 15459
rect 10439 15069 10473 15117
rect 11649 15069 11683 15117
rect 11915 14971 11949 15099
rect 13125 14971 13159 15099
rect 10469 14667 10503 14835
rect 11679 14667 11713 14835
rect 11915 14611 11949 14739
rect 13125 14611 13159 14739
rect 10469 14243 10503 14411
rect 11679 14243 11713 14411
rect 11915 14251 11949 14379
rect 13125 14251 13159 14379
rect 5858 13665 5892 13793
rect 7068 13665 7102 13793
rect 7334 13701 7368 13749
rect 8544 13701 8578 13749
rect 5858 13305 5892 13433
rect 7068 13305 7102 13433
rect 7334 13403 7368 13451
rect 8544 13403 8578 13451
rect 5858 12945 5892 13073
rect 7068 12945 7102 13073
rect 7304 13001 7338 13169
rect 8514 13001 8548 13169
rect 5858 12585 5892 12713
rect 7068 12585 7102 12713
rect 7304 12577 7338 12745
rect 8514 12577 8548 12745
rect 8982 13696 9016 13824
rect 9310 13696 9344 13824
rect 8982 13288 9016 13416
rect 9310 13288 9344 13416
rect 8982 12602 9016 12970
rect 9310 12602 9344 12970
rect 9673 13696 9707 13824
rect 10001 13696 10035 13824
rect 9673 13288 9707 13416
rect 10001 13288 10035 13416
rect 9673 12602 9707 12970
rect 10001 12602 10035 12970
rect 10439 13701 10473 13749
rect 11649 13701 11683 13749
rect 11915 13665 11949 13793
rect 13125 13665 13159 13793
rect 10439 13403 10473 13451
rect 11649 13403 11683 13451
rect 11915 13305 11949 13433
rect 13125 13305 13159 13433
rect 10469 13001 10503 13169
rect 11679 13001 11713 13169
rect 11915 12945 11949 13073
rect 13125 12945 13159 13073
rect 10469 12577 10503 12745
rect 11679 12577 11713 12745
rect 11915 12585 11949 12713
rect 13125 12585 13159 12713
rect 5858 11999 5892 12127
rect 7068 11999 7102 12127
rect 7334 12035 7368 12083
rect 8544 12035 8578 12083
rect 5858 11639 5892 11767
rect 7068 11639 7102 11767
rect 7334 11737 7368 11785
rect 8544 11737 8578 11785
rect 5858 11279 5892 11407
rect 7068 11279 7102 11407
rect 7304 11335 7338 11503
rect 8514 11335 8548 11503
rect 5858 10919 5892 11047
rect 7068 10919 7102 11047
rect 7304 10911 7338 11079
rect 8514 10911 8548 11079
rect 8982 12030 9016 12158
rect 9310 12030 9344 12158
rect 8982 11622 9016 11750
rect 9310 11622 9344 11750
rect 8982 10936 9016 11304
rect 9310 10936 9344 11304
rect 9673 12030 9707 12158
rect 10001 12030 10035 12158
rect 9673 11622 9707 11750
rect 10001 11622 10035 11750
rect 9673 10936 9707 11304
rect 10001 10936 10035 11304
rect 10439 12035 10473 12083
rect 11649 12035 11683 12083
rect 11915 11999 11949 12127
rect 13125 11999 13159 12127
rect 10439 11737 10473 11785
rect 11649 11737 11683 11785
rect 11915 11639 11949 11767
rect 13125 11639 13159 11767
rect 10469 11335 10503 11503
rect 11679 11335 11713 11503
rect 11915 11279 11949 11407
rect 13125 11279 13159 11407
rect 10469 10911 10503 11079
rect 11679 10911 11713 11079
rect 11915 10919 11949 11047
rect 13125 10919 13159 11047
rect 5858 10333 5892 10461
rect 7068 10333 7102 10461
rect 7334 10369 7368 10417
rect 8544 10369 8578 10417
rect 5858 9973 5892 10101
rect 7068 9973 7102 10101
rect 7334 10071 7368 10119
rect 8544 10071 8578 10119
rect 5858 9613 5892 9741
rect 7068 9613 7102 9741
rect 7304 9669 7338 9837
rect 8514 9669 8548 9837
rect 5858 9253 5892 9381
rect 7068 9253 7102 9381
rect 7304 9245 7338 9413
rect 8514 9245 8548 9413
rect 8982 10364 9016 10492
rect 9310 10364 9344 10492
rect 8982 9956 9016 10084
rect 9310 9956 9344 10084
rect 8982 9270 9016 9638
rect 9310 9270 9344 9638
rect 9673 10364 9707 10492
rect 10001 10364 10035 10492
rect 9673 9956 9707 10084
rect 10001 9956 10035 10084
rect 9673 9270 9707 9638
rect 10001 9270 10035 9638
rect 10439 10369 10473 10417
rect 11649 10369 11683 10417
rect 11915 10333 11949 10461
rect 13125 10333 13159 10461
rect 10439 10071 10473 10119
rect 11649 10071 11683 10119
rect 11915 9973 11949 10101
rect 13125 9973 13159 10101
rect 10469 9669 10503 9837
rect 11679 9669 11713 9837
rect 11915 9613 11949 9741
rect 13125 9613 13159 9741
rect 10469 9245 10503 9413
rect 11679 9245 11713 9413
rect 11915 9253 11949 9381
rect 13125 9253 13159 9381
rect 5858 8667 5892 8795
rect 7068 8667 7102 8795
rect 7334 8703 7368 8751
rect 8544 8703 8578 8751
rect 5858 8307 5892 8435
rect 7068 8307 7102 8435
rect 7334 8405 7368 8453
rect 8544 8405 8578 8453
rect 5858 7947 5892 8075
rect 7068 7947 7102 8075
rect 7304 8003 7338 8171
rect 8514 8003 8548 8171
rect 5858 7587 5892 7715
rect 7068 7587 7102 7715
rect 7304 7579 7338 7747
rect 8514 7579 8548 7747
rect 8982 8698 9016 8826
rect 9310 8698 9344 8826
rect 8982 8290 9016 8418
rect 9310 8290 9344 8418
rect 8982 7604 9016 7972
rect 9310 7604 9344 7972
rect 9673 8698 9707 8826
rect 10001 8698 10035 8826
rect 9673 8290 9707 8418
rect 10001 8290 10035 8418
rect 9673 7604 9707 7972
rect 10001 7604 10035 7972
rect 10439 8703 10473 8751
rect 11649 8703 11683 8751
rect 11915 8667 11949 8795
rect 13125 8667 13159 8795
rect 10439 8405 10473 8453
rect 11649 8405 11683 8453
rect 11915 8307 11949 8435
rect 13125 8307 13159 8435
rect 10469 8003 10503 8171
rect 11679 8003 11713 8171
rect 11915 7947 11949 8075
rect 13125 7947 13159 8075
rect 10469 7579 10503 7747
rect 11679 7579 11713 7747
rect 11915 7587 11949 7715
rect 13125 7587 13159 7715
rect 15117 17732 15155 17766
rect 15117 15884 15155 15918
rect 16166 17288 16200 17434
rect 17476 17288 17510 17434
rect 16166 16918 16200 17064
rect 17476 16918 17510 17064
rect 16548 16694 17136 16728
rect 17436 16622 17614 16656
rect 17436 16348 17614 16382
rect 16548 16240 17136 16274
rect 14901 12694 14935 13440
rect 15207 12694 15241 13440
rect 15401 12694 15435 13440
rect 15707 12694 15741 13440
rect 15901 12694 15935 13440
rect 16207 12694 16241 13440
rect 16401 12694 16435 13440
rect 16707 12694 16741 13440
rect 16901 12694 16935 13440
rect 17207 12694 17241 13440
rect 17401 12694 17435 13440
rect 17707 12694 17741 13440
rect 14564 11712 14818 11746
rect 14564 10564 14818 10598
rect 14564 10456 14818 10490
rect 14564 9308 14818 9342
rect 17005 11243 17039 11285
rect 18167 11243 18201 11285
rect 16948 9996 16982 10218
rect 18290 9996 18324 10218
rect 16948 9396 16982 9618
rect 18290 9396 18324 9618
rect 14538 8636 14638 8670
rect 14938 8636 15038 8670
rect 15338 8636 15438 8670
rect 15738 8636 15838 8670
rect 16138 8636 16238 8670
rect 16538 8636 16638 8670
rect 16938 8636 17038 8670
rect 17338 8636 17438 8670
rect 17738 8636 17838 8670
rect 18138 8636 18238 8670
rect 14538 7506 14638 7540
rect 14938 7506 15038 7540
rect 15338 7506 15438 7540
rect 15738 7506 15838 7540
rect 16138 7506 16238 7540
rect 16538 7506 16638 7540
rect 16938 7506 17038 7540
rect 17338 7506 17438 7540
rect 17738 7506 17838 7540
rect 18138 7506 18238 7540
<< locali >>
rect -1047 19784 18654 20384
rect -1047 19683 764 19784
rect 5507 19732 12606 19784
rect 5460 19716 12672 19732
rect -1047 19530 -564 19683
rect 4357 19613 4673 19683
rect 4357 19530 4507 19613
rect -1047 19401 784 19530
rect -1047 7535 -560 19401
rect -436 19198 784 19401
rect 1061 19445 2822 19453
rect 1061 19413 4304 19445
rect 1061 19397 2943 19413
rect -436 19110 -99 19198
rect 576 19110 784 19198
rect -436 19100 -85 19110
rect -436 18723 -269 19100
rect -436 15674 -269 15811
rect -200 19029 -85 19100
rect 423 19029 495 19110
rect -200 18995 -69 19029
rect 407 18995 495 19029
rect -200 18967 -85 18995
rect -200 18799 -153 18967
rect -119 18799 -85 18967
rect -200 18771 -85 18799
rect 423 18967 495 18995
rect 423 18799 457 18967
rect 491 18799 495 18967
rect 423 18771 495 18799
rect -200 18737 -69 18771
rect 407 18737 495 18771
rect -200 18702 495 18737
rect 582 19035 784 19110
rect -85 18579 -69 18613
rect 407 18579 423 18613
rect -153 18551 -119 18567
rect -153 18367 -119 18383
rect 457 18551 527 18567
rect 491 18383 527 18551
rect 457 18367 527 18383
rect -85 18321 -69 18355
rect 407 18321 423 18355
rect -200 18286 423 18321
rect -85 18163 -69 18197
rect 407 18163 423 18197
rect 491 18151 527 18367
rect -153 18135 -119 18151
rect -153 17951 -119 17967
rect 457 18135 527 18151
rect 491 17967 527 18135
rect 457 17951 527 17967
rect -85 17905 -69 17939
rect 407 17905 423 17939
rect -200 17870 423 17905
rect -85 17747 -69 17781
rect 407 17747 423 17781
rect 491 17735 527 17951
rect -153 17719 -119 17735
rect -153 17535 -119 17551
rect 457 17719 527 17735
rect 491 17551 527 17719
rect 457 17535 527 17551
rect -85 17489 -69 17523
rect 407 17489 423 17523
rect -200 17454 423 17489
rect -85 17331 -69 17365
rect 407 17331 423 17365
rect 491 17319 527 17535
rect -153 17303 -119 17319
rect -153 17119 -119 17135
rect 457 17303 527 17319
rect 491 17135 527 17303
rect 457 17119 527 17135
rect -85 17073 -69 17107
rect 407 17073 423 17107
rect -200 17038 423 17073
rect -85 16915 -69 16949
rect 407 16915 423 16949
rect 491 16903 527 17119
rect -153 16887 -119 16903
rect -153 16703 -119 16719
rect 457 16887 527 16903
rect 491 16719 527 16887
rect 457 16703 527 16719
rect -85 16657 -69 16691
rect 407 16657 423 16691
rect -200 16622 423 16657
rect -85 16499 -69 16533
rect 407 16499 423 16533
rect 491 16487 527 16703
rect -153 16471 -119 16487
rect -153 16287 -119 16303
rect 457 16471 527 16487
rect 491 16303 527 16471
rect 457 16287 527 16303
rect -85 16241 -69 16275
rect 407 16241 423 16275
rect -200 16206 423 16241
rect -157 16083 -69 16117
rect 407 16083 495 16117
rect -157 16055 -85 16083
rect -157 15887 -153 16055
rect -119 15887 -85 16055
rect -157 15859 -85 15887
rect 423 16055 495 16083
rect 423 15887 457 16055
rect 491 15887 495 16055
rect 423 15859 495 15887
rect -157 15825 -69 15859
rect 407 15825 495 15859
rect -200 15790 495 15825
rect -200 15702 -85 15790
rect 423 15702 495 15790
rect 633 15793 784 19035
rect 582 15702 784 15793
rect -200 15674 -115 15702
rect -436 15621 -115 15674
rect -157 15614 -115 15621
rect 560 15614 784 15702
rect 332 14846 784 15614
rect 1057 19363 1117 19397
rect 2631 19379 2943 19397
rect 4314 19379 4374 19413
rect 2631 19363 4374 19379
rect 1057 19353 4374 19363
rect 1057 19337 2883 19353
rect 1091 19325 2657 19337
rect 1340 19279 1832 19325
rect 1340 19245 1402 19279
rect 1770 19245 1832 19279
rect 1340 19186 1386 19245
rect 1374 19110 1386 19186
rect 1340 19051 1386 19110
rect 1786 19186 1832 19245
rect 1786 19110 1798 19186
rect 1786 19051 1832 19110
rect 1340 19017 1402 19051
rect 1770 19017 1832 19051
rect 2040 19279 2532 19325
rect 2040 19245 2102 19279
rect 2470 19245 2532 19279
rect 2040 19186 2086 19245
rect 2074 19110 2086 19186
rect 2040 19051 2086 19110
rect 2486 19186 2532 19245
rect 2486 19110 2498 19186
rect 2486 19051 2532 19110
rect 2040 19017 2102 19051
rect 2470 19017 2532 19051
rect 1260 18861 1402 18895
rect 1770 18861 1786 18895
rect 2086 18861 2102 18895
rect 2470 18861 2486 18895
rect 1260 18267 1294 18861
rect 1340 18802 1374 18818
rect 1340 18310 1374 18326
rect 1798 18802 1832 18818
rect 2040 18802 2074 18818
rect 1832 18603 2040 18624
rect 1832 18539 1898 18603
rect 1954 18539 2040 18603
rect 1832 18517 2040 18539
rect 1798 18310 1832 18326
rect 2040 18310 2074 18326
rect 2498 18802 2532 18818
rect 2532 18509 2657 18634
rect 2498 18310 2532 18326
rect 1260 18233 1402 18267
rect 1770 18233 1786 18267
rect 2086 18233 2102 18267
rect 2470 18233 2486 18267
rect 1386 18077 1402 18111
rect 1770 18077 1786 18111
rect 2086 18077 2102 18111
rect 2470 18077 2486 18111
rect 1340 18018 1374 18034
rect 1340 17526 1374 17542
rect 1798 18018 1832 18034
rect 2040 18018 2074 18034
rect 1832 17716 2040 17823
rect 1798 17526 1832 17542
rect 1386 17449 1402 17483
rect 1770 17449 1786 17483
rect 1386 17293 1402 17327
rect 1770 17293 1786 17327
rect 1340 17234 1374 17250
rect 1340 16742 1374 16758
rect 1798 17234 1832 17250
rect 1876 17049 1972 17716
rect 2040 17526 2074 17542
rect 2498 18018 2532 18034
rect 2532 17719 2657 17844
rect 2498 17526 2532 17542
rect 2086 17449 2102 17483
rect 2470 17449 2486 17483
rect 2086 17293 2102 17327
rect 2470 17293 2486 17327
rect 2040 17234 2074 17250
rect 1832 16942 2040 17049
rect 1798 16742 1832 16758
rect 2040 16742 2074 16758
rect 2498 17234 2532 17250
rect 2532 16935 2657 17060
rect 2498 16742 2532 16758
rect 1386 16665 1402 16699
rect 1770 16665 1786 16699
rect 2086 16665 2102 16699
rect 2470 16665 2486 16699
rect 1244 16509 1402 16543
rect 1770 16509 1786 16543
rect 2086 16509 2102 16543
rect 2470 16509 2486 16543
rect 1244 15964 1278 16509
rect 1149 15945 1278 15964
rect 1340 16450 1374 16466
rect 1340 15958 1374 15974
rect 1798 16450 1832 16466
rect 2040 16450 2074 16466
rect 1832 16241 2040 16263
rect 1832 16177 1901 16241
rect 1957 16177 2040 16241
rect 1832 16156 2040 16177
rect 1798 15958 1832 15974
rect 2040 15958 2074 15974
rect 2498 16450 2532 16466
rect 2532 16143 2657 16268
rect 2498 15958 2532 15974
rect 1149 15765 1167 15945
rect 1256 15915 1278 15945
rect 1256 15881 1402 15915
rect 1770 15881 1786 15915
rect 2086 15881 2102 15915
rect 2470 15881 2486 15915
rect 1256 15765 1278 15881
rect 1149 15735 1278 15765
rect 1057 15437 1091 15453
rect 1340 15725 1402 15759
rect 1770 15725 1832 15759
rect 1340 15666 1386 15725
rect 1374 15590 1386 15666
rect 1340 15531 1386 15590
rect 1786 15666 1832 15725
rect 1786 15590 1798 15666
rect 1786 15531 1832 15590
rect 1340 15497 1402 15531
rect 1770 15497 1832 15531
rect 1340 15437 1832 15497
rect 2040 15725 2102 15759
rect 2470 15725 2532 15759
rect 2040 15666 2086 15725
rect 2074 15590 2086 15666
rect 2040 15531 2086 15590
rect 2486 15666 2532 15725
rect 2486 15590 2498 15666
rect 2486 15531 2532 15590
rect 2040 15497 2102 15531
rect 2470 15497 2532 15531
rect 2040 15437 2532 15497
rect 2691 15453 2883 19337
rect 2657 15437 2883 15453
rect 1057 15427 2883 15437
rect 1057 15393 1117 15427
rect 2631 15393 2883 15427
rect 1073 15334 2883 15393
rect -436 14773 -4 14846
rect 2394 14773 2549 14846
rect -436 14754 1 14773
rect -436 14079 -203 14754
rect -115 14689 1 14754
rect 2358 14770 2549 14773
rect 2358 14689 2461 14770
rect -115 14685 300 14689
rect 2053 14685 2461 14689
rect -115 14651 70 14685
rect 238 14651 300 14685
rect 470 14651 486 14685
rect 654 14651 670 14685
rect 886 14651 902 14685
rect 1070 14651 1086 14685
rect 1302 14651 1318 14685
rect 1486 14651 1502 14685
rect 1718 14651 1734 14685
rect 1902 14651 1918 14685
rect 2053 14651 2150 14685
rect 2318 14651 2461 14685
rect -115 14617 300 14651
rect 2053 14617 2461 14651
rect -115 14601 42 14617
rect -115 14125 8 14601
rect -115 14109 42 14125
rect 266 14601 300 14617
rect 266 14109 300 14125
rect -115 14079 300 14109
rect -436 14075 300 14079
rect -436 14041 70 14075
rect 238 14041 300 14075
rect -436 14037 300 14041
rect 389 14601 458 14617
rect 389 14125 424 14601
rect 389 14109 458 14125
rect 682 14601 716 14617
rect 682 14109 716 14125
rect 805 14601 874 14617
rect 805 14125 840 14601
rect 805 14109 874 14125
rect 1098 14601 1132 14617
rect 1098 14109 1132 14125
rect 1221 14601 1290 14617
rect 1221 14125 1256 14601
rect 1221 14109 1290 14125
rect 1514 14601 1548 14617
rect 1514 14109 1548 14125
rect 1637 14601 1706 14617
rect 1637 14125 1672 14601
rect 1637 14109 1706 14125
rect 1930 14601 1964 14617
rect 1930 14109 1964 14125
rect 2053 14601 2122 14617
rect 2053 14125 2088 14601
rect 2053 14109 2122 14125
rect 2346 14601 2461 14617
rect 2380 14125 2461 14601
rect 2346 14109 2461 14125
rect -436 13903 -115 14037
rect -27 13999 8 14037
rect 389 13903 424 14109
rect 470 14041 486 14075
rect 654 14041 670 14075
rect 805 13992 840 14109
rect 886 14041 902 14075
rect 1070 14041 1086 14075
rect 1221 14004 1256 14109
rect 1302 14041 1318 14075
rect 1486 14041 1502 14075
rect 1221 13992 1257 14004
rect 805 13983 1257 13992
rect 805 13954 964 13983
rect 941 13946 964 13954
rect 1084 13954 1257 13983
rect 1084 13946 1114 13954
rect 941 13939 1114 13946
rect 1637 13903 1672 14109
rect 2053 14095 2461 14109
rect 2549 14095 2550 14109
rect 2053 14075 2550 14095
rect 1718 14041 1734 14075
rect 1902 14041 1918 14075
rect 2053 14041 2150 14075
rect 2318 14041 2550 14075
rect 2053 14037 2550 14041
rect 2053 13999 2088 14037
rect 2358 13905 2551 14037
rect 1881 13903 1897 13905
rect -436 13836 -213 13903
rect -229 13809 -213 13836
rect 393 13869 595 13903
rect 1723 13869 1897 13903
rect 393 13854 533 13869
rect 393 13809 409 13854
rect 499 13807 533 13854
rect 1785 13829 1897 13869
rect 2527 13829 2551 13905
rect 1785 13807 1819 13829
rect 659 13767 675 13801
rect 1643 13767 1659 13801
rect 613 13717 647 13733
rect 533 13575 613 13676
rect 613 13525 647 13541
rect 1671 13717 1705 13733
rect 1671 13525 1705 13541
rect 659 13457 675 13491
rect 1643 13457 1659 13491
rect 499 13389 533 13451
rect 1785 13389 1819 13451
rect 499 13355 595 13389
rect 1723 13355 1819 13389
rect 1154 13218 1398 13251
rect 1154 13005 1185 13218
rect 1366 13005 1398 13218
rect 1154 12960 1398 13005
rect 1190 12840 1365 12960
rect 2467 12860 2584 12876
rect -346 12806 -250 12840
rect 2232 12806 2328 12840
rect -346 12744 -312 12806
rect -167 12726 241 12806
rect -167 12692 -151 12726
rect 225 12692 241 12726
rect 469 12726 877 12806
rect 469 12692 485 12726
rect 861 12692 877 12726
rect 1105 12726 1513 12806
rect 1105 12692 1121 12726
rect 1497 12692 1513 12726
rect 1741 12726 2149 12806
rect 1741 12692 1757 12726
rect 2133 12692 2149 12726
rect 2294 12744 2328 12806
rect -244 12664 -210 12680
rect -244 12580 -210 12596
rect 284 12664 318 12680
rect 284 12580 318 12596
rect 392 12664 426 12680
rect 392 12580 426 12596
rect 920 12664 954 12680
rect 920 12580 954 12596
rect 1028 12664 1062 12680
rect 1028 12580 1062 12596
rect 1556 12664 1590 12680
rect 1556 12580 1590 12596
rect 1664 12664 1698 12680
rect 1664 12580 1698 12596
rect 2192 12664 2226 12680
rect 2192 12580 2226 12596
rect -167 12534 -151 12568
rect 225 12534 241 12568
rect 469 12534 485 12568
rect 861 12534 877 12568
rect 1105 12534 1121 12568
rect 1497 12534 1513 12568
rect 1741 12534 1757 12568
rect 2133 12534 2149 12568
rect -346 12454 -312 12516
rect 2294 12454 2328 12516
rect -346 12420 -250 12454
rect 2232 12420 2328 12454
rect 44 12409 166 12420
rect 44 12308 62 12409
rect 146 12308 166 12409
rect 2184 12353 2467 12356
rect 44 12281 166 12308
rect 2059 12331 2467 12353
rect 2059 12294 2207 12331
rect 298 12179 314 12294
rect 2111 12260 2207 12294
rect 2111 12179 2467 12260
rect 320 12009 438 12179
rect 2059 12166 2467 12179
rect -436 11649 438 12009
rect 619 12048 715 12082
rect 2237 12048 2333 12082
rect 619 11986 653 12048
rect 749 11986 2333 12048
rect 749 11980 2299 11986
rect 749 11972 795 11980
rect 779 11946 795 11972
rect 2157 11946 2299 11980
rect 733 11887 767 11903
rect 733 11719 767 11735
rect 2185 11887 2299 11946
rect 2219 11735 2299 11887
rect 2185 11676 2299 11735
rect 779 11651 795 11676
rect 619 11574 653 11636
rect 751 11642 795 11651
rect 2157 11642 2299 11676
rect 751 11636 2299 11642
rect 751 11574 2333 11636
rect 619 11540 715 11574
rect 2237 11540 2333 11574
rect 666 11510 925 11540
rect 666 11357 698 11510
rect 875 11357 925 11510
rect 666 11315 925 11357
rect 241 11170 301 11204
rect 2297 11170 2357 11204
rect 241 11144 275 11170
rect 2237 11144 2357 11170
rect 401 11078 1117 11101
rect 401 11044 417 11078
rect 939 11061 1117 11078
rect 939 11044 955 11061
rect 355 10985 389 11001
rect 355 10307 389 10323
rect 967 10985 1001 11001
rect 967 10307 1001 10323
rect 401 10230 417 10264
rect 939 10237 955 10264
rect 1076 10237 1117 11061
rect 1395 11038 1411 11072
rect 2179 11038 2195 11072
rect 2237 10995 2323 11144
rect 1349 10979 1383 10995
rect 1349 10887 1383 10903
rect 2207 10979 2323 10995
rect 2241 10903 2323 10979
rect 2207 10887 2323 10903
rect 1395 10810 1411 10844
rect 2179 10810 2195 10844
rect 1321 10646 1337 10680
rect 2181 10646 2197 10680
rect 2237 10603 2323 10887
rect 1275 10587 1309 10603
rect 939 10230 1275 10237
rect 401 10198 1275 10230
rect 1275 10121 1309 10137
rect 2209 10587 2323 10603
rect 2243 10137 2323 10587
rect 2209 10121 2323 10137
rect 1321 10044 1337 10078
rect 2181 10044 2197 10078
rect 241 9943 275 9969
rect 2237 9969 2323 10121
rect 2237 9943 2357 9969
rect 241 9909 301 9943
rect 2297 9909 2357 9943
rect 1253 9521 2351 9909
rect 2584 12166 2589 12353
rect 2467 9756 2584 9772
rect 2802 9521 2883 15334
rect 1253 9425 2883 9521
rect 973 9391 1033 9425
rect 2373 9391 2883 9425
rect 973 9365 1007 9391
rect 2399 9365 2883 9391
rect 1155 9299 1171 9333
rect 1539 9299 1555 9333
rect 1855 9299 1871 9333
rect 2239 9299 2255 9333
rect 1109 9240 1143 9256
rect 1109 8748 1143 8764
rect 1567 9240 1601 9256
rect 1567 8748 1601 8764
rect 1809 9240 1843 9256
rect 1809 8748 1843 8764
rect 2267 9240 2399 9256
rect 2301 8764 2399 9240
rect 2433 9116 2883 9365
rect 2267 8748 2399 8764
rect 1155 8671 1171 8705
rect 1539 8671 1555 8705
rect 1855 8671 1871 8705
rect 2239 8671 2255 8705
rect 1155 8515 1171 8549
rect 1539 8515 1555 8549
rect 1855 8515 1871 8549
rect 2239 8515 2255 8549
rect 2301 8472 2399 8748
rect 2762 8504 2883 9116
rect 1109 8456 1143 8472
rect 1109 7964 1143 7980
rect 1567 8456 1601 8472
rect 1567 7964 1601 7980
rect 1809 8456 1843 8472
rect 1809 7964 1843 7980
rect 2267 8456 2399 8472
rect 2301 7980 2399 8456
rect 2267 7964 2399 7980
rect 1155 7887 1171 7921
rect 1539 7887 1555 7921
rect 1855 7887 1871 7921
rect 2239 7887 2255 7921
rect 973 7817 1007 7843
rect 2433 8403 2883 8504
rect 2399 7817 2433 7843
rect 973 7783 1033 7817
rect 2373 7783 2433 7817
rect 2651 7638 2883 8403
rect 2917 19295 4340 19353
rect 2917 19277 3098 19295
rect 3036 19261 3098 19277
rect 3466 19277 3798 19295
rect 3466 19261 3528 19277
rect 3036 19218 3082 19261
rect 3482 19218 3528 19261
rect 3036 19202 3070 19218
rect 3036 19110 3070 19126
rect 3494 19202 3528 19218
rect 3494 19110 3528 19126
rect 3736 19261 3798 19277
rect 4166 19261 4340 19295
rect 3736 19218 3782 19261
rect 4182 19218 4340 19261
rect 3736 19202 3770 19218
rect 3736 19110 3770 19126
rect 4194 19202 4340 19218
rect 4228 19126 4340 19202
rect 4194 19110 4340 19126
rect 3082 19033 3098 19067
rect 3466 19033 3482 19067
rect 3782 19033 3798 19067
rect 4166 19033 4182 19067
rect 3082 18877 3098 18911
rect 3466 18877 3482 18911
rect 3782 18877 3798 18911
rect 4166 18877 4182 18911
rect 4216 18834 4340 19110
rect 3036 18818 3070 18834
rect 3036 18326 3070 18342
rect 3494 18818 3528 18834
rect 3494 18326 3528 18342
rect 3736 18818 3770 18834
rect 3736 18326 3770 18342
rect 4194 18818 4340 18834
rect 4228 18342 4340 18818
rect 4194 18326 4340 18342
rect 3082 18249 3098 18283
rect 3466 18249 3482 18283
rect 3782 18249 3798 18283
rect 4166 18249 4182 18283
rect 3082 18093 3098 18127
rect 3466 18093 3482 18127
rect 3782 18093 3798 18127
rect 4166 18093 4182 18127
rect 4216 18050 4340 18326
rect 3036 18034 3070 18050
rect 3036 17542 3070 17558
rect 3494 18034 3528 18050
rect 3494 17542 3528 17558
rect 3736 18034 3770 18050
rect 3736 17542 3770 17558
rect 4194 18034 4340 18050
rect 4228 17558 4340 18034
rect 4194 17542 4340 17558
rect 3082 17465 3098 17499
rect 3466 17465 3482 17499
rect 3782 17465 3798 17499
rect 4166 17465 4182 17499
rect 3082 17309 3098 17343
rect 3466 17309 3482 17343
rect 3782 17309 3798 17343
rect 4166 17309 4182 17343
rect 4216 17266 4340 17542
rect 3036 17250 3070 17266
rect 3036 16758 3070 16774
rect 3494 17250 3528 17266
rect 3494 16758 3528 16774
rect 3736 17250 3770 17266
rect 3736 16758 3770 16774
rect 4194 17250 4340 17266
rect 4228 16774 4340 17250
rect 4194 16758 4340 16774
rect 3082 16681 3098 16715
rect 3466 16681 3482 16715
rect 3782 16681 3798 16715
rect 4166 16681 4182 16715
rect 3082 16525 3098 16559
rect 3466 16525 3482 16559
rect 3782 16525 3798 16559
rect 4166 16525 4182 16559
rect 4216 16482 4340 16758
rect 3036 16466 3070 16482
rect 3036 15974 3070 15990
rect 3494 16466 3528 16482
rect 3494 15974 3528 15990
rect 3736 16466 3770 16482
rect 3736 15974 3770 15990
rect 4194 16466 4340 16482
rect 4228 15990 4340 16466
rect 4194 15974 4340 15990
rect 3082 15897 3098 15931
rect 3466 15897 3482 15931
rect 3782 15897 3798 15931
rect 4166 15897 4182 15931
rect 3082 15741 3098 15775
rect 3466 15741 3482 15775
rect 3782 15741 3798 15775
rect 4166 15741 4182 15775
rect 4216 15698 4340 15974
rect 3036 15682 3070 15698
rect 3036 15190 3070 15206
rect 3494 15682 3528 15698
rect 3494 15190 3528 15206
rect 3736 15682 3770 15698
rect 3736 15190 3770 15206
rect 4194 15682 4340 15698
rect 4228 15206 4340 15682
rect 4194 15190 4340 15206
rect 3082 15113 3098 15147
rect 3466 15113 3482 15147
rect 3782 15113 3798 15147
rect 4166 15113 4182 15147
rect 3082 14957 3098 14991
rect 3466 14957 3482 14991
rect 3782 14957 3798 14991
rect 4166 14957 4182 14991
rect 4216 14914 4340 15190
rect 3036 14898 3070 14914
rect 3036 14406 3070 14422
rect 3494 14898 3528 14914
rect 3736 14898 3770 14914
rect 3528 14699 3736 14720
rect 3528 14635 3594 14699
rect 3650 14635 3736 14699
rect 3528 14613 3736 14635
rect 3494 14406 3528 14422
rect 3736 14406 3770 14422
rect 4194 14898 4340 14914
rect 4228 14422 4340 14898
rect 4194 14406 4340 14422
rect 3082 14329 3098 14363
rect 3466 14329 3482 14363
rect 3782 14329 3798 14363
rect 4166 14329 4182 14363
rect 3082 14173 3098 14207
rect 3466 14173 3482 14207
rect 3782 14173 3798 14207
rect 4166 14173 4182 14207
rect 4216 14130 4340 14406
rect 3036 14114 3070 14130
rect 3036 13622 3070 13638
rect 3494 14114 3528 14130
rect 3736 14114 3770 14130
rect 3528 13812 3736 13919
rect 3494 13622 3528 13638
rect 3082 13545 3098 13579
rect 3466 13545 3482 13579
rect 3082 13389 3098 13423
rect 3466 13389 3482 13423
rect 3036 13330 3070 13346
rect 3036 12838 3070 12854
rect 3494 13330 3528 13346
rect 3572 13145 3668 13812
rect 3736 13622 3770 13638
rect 4194 14114 4340 14130
rect 4228 13638 4340 14114
rect 4194 13622 4340 13638
rect 3782 13545 3798 13579
rect 4166 13545 4182 13579
rect 3782 13389 3798 13423
rect 4166 13389 4182 13423
rect 4216 13346 4340 13622
rect 3736 13330 3770 13346
rect 3528 13038 3736 13145
rect 3494 12838 3528 12854
rect 3736 12838 3770 12854
rect 4194 13330 4340 13346
rect 4228 12854 4340 13330
rect 4194 12838 4340 12854
rect 3082 12761 3098 12795
rect 3466 12761 3482 12795
rect 3782 12761 3798 12795
rect 4166 12761 4182 12795
rect 3082 12605 3098 12639
rect 3466 12605 3482 12639
rect 3782 12605 3798 12639
rect 4166 12605 4182 12639
rect 4216 12562 4340 12838
rect 3036 12546 3070 12562
rect 3036 12054 3070 12070
rect 3494 12546 3528 12562
rect 3736 12546 3770 12562
rect 3528 12337 3736 12359
rect 3528 12273 3597 12337
rect 3653 12273 3736 12337
rect 3528 12252 3736 12273
rect 3494 12054 3528 12070
rect 3736 12054 3770 12070
rect 4194 12546 4340 12562
rect 4228 12070 4340 12546
rect 4194 12054 4340 12070
rect 3082 11977 3098 12011
rect 3466 11977 3482 12011
rect 3782 11977 3798 12011
rect 4166 11977 4182 12011
rect 3082 11821 3098 11855
rect 3466 11821 3482 11855
rect 3782 11821 3798 11855
rect 4166 11821 4182 11855
rect 4216 11778 4340 12054
rect 3036 11762 3070 11778
rect 3036 11270 3070 11286
rect 3494 11762 3528 11778
rect 3494 11270 3528 11286
rect 3736 11762 3770 11778
rect 3736 11270 3770 11286
rect 4194 11762 4340 11778
rect 4228 11286 4340 11762
rect 4194 11270 4340 11286
rect 3082 11193 3098 11227
rect 3466 11193 3482 11227
rect 3782 11193 3798 11227
rect 4166 11193 4182 11227
rect 3082 11037 3098 11071
rect 3466 11037 3482 11071
rect 3782 11037 3798 11071
rect 4166 11037 4182 11071
rect 4216 10994 4340 11270
rect 3036 10978 3070 10994
rect 3036 10486 3070 10502
rect 3494 10978 3528 10994
rect 3494 10486 3528 10502
rect 3736 10978 3770 10994
rect 3736 10486 3770 10502
rect 4194 10978 4340 10994
rect 4228 10502 4340 10978
rect 4194 10486 4340 10502
rect 3082 10409 3098 10443
rect 3466 10409 3482 10443
rect 3782 10409 3798 10443
rect 4166 10409 4182 10443
rect 3082 10253 3098 10287
rect 3466 10253 3482 10287
rect 3782 10253 3798 10287
rect 4166 10253 4182 10287
rect 4216 10210 4340 10486
rect 3036 10194 3070 10210
rect 3036 9702 3070 9718
rect 3494 10194 3528 10210
rect 3494 9702 3528 9718
rect 3736 10194 3770 10210
rect 3736 9702 3770 9718
rect 4194 10194 4340 10210
rect 4228 9718 4340 10194
rect 4194 9702 4340 9718
rect 3082 9625 3098 9659
rect 3466 9625 3482 9659
rect 3782 9625 3798 9659
rect 4166 9625 4182 9659
rect 3082 9469 3098 9503
rect 3466 9469 3482 9503
rect 3782 9469 3798 9503
rect 4166 9469 4182 9503
rect 4216 9426 4340 9702
rect 3036 9410 3070 9426
rect 3036 8918 3070 8934
rect 3494 9410 3528 9426
rect 3494 8918 3528 8934
rect 3736 9410 3770 9426
rect 3736 8918 3770 8934
rect 4194 9410 4340 9426
rect 4228 8934 4340 9410
rect 4194 8918 4340 8934
rect 3082 8841 3098 8875
rect 3466 8841 3482 8875
rect 3782 8841 3798 8875
rect 4166 8841 4182 8875
rect 3082 8685 3098 8719
rect 3466 8685 3482 8719
rect 3782 8685 3798 8719
rect 4166 8685 4182 8719
rect 4216 8642 4340 8918
rect 3036 8626 3070 8642
rect 3036 8134 3070 8150
rect 3494 8626 3528 8642
rect 3494 8134 3528 8150
rect 3736 8626 3770 8642
rect 3736 8134 3770 8150
rect 4194 8626 4340 8642
rect 4228 8150 4340 8626
rect 4194 8134 4340 8150
rect 3082 8057 3098 8091
rect 3466 8057 3482 8091
rect 3782 8057 3798 8091
rect 4166 8057 4182 8091
rect 3082 7901 3098 7935
rect 3466 7901 3482 7935
rect 3782 7901 3798 7935
rect 4166 7901 4182 7935
rect 4216 7858 4340 8134
rect 3036 7846 3070 7858
rect 2917 7842 3070 7846
rect 2917 7766 3036 7842
rect 2917 7750 3070 7766
rect 3494 7842 3528 7858
rect 3494 7750 3528 7766
rect 2917 7707 3082 7750
rect 3482 7707 3528 7750
rect 2917 7673 3098 7707
rect 3466 7678 3528 7707
rect 3736 7842 3770 7858
rect 3736 7750 3770 7766
rect 4194 7842 4340 7858
rect 4228 7766 4340 7842
rect 4194 7750 4340 7766
rect 3736 7707 3782 7750
rect 4182 7707 4340 7750
rect 3736 7678 3798 7707
rect 3466 7673 3798 7678
rect 4166 7673 4340 7707
rect 2917 7638 4340 7673
rect 2651 7612 4374 7638
rect 2651 7591 2943 7612
rect 2883 7578 2943 7591
rect 4314 7578 4374 7612
rect -1047 7379 -436 7535
rect -1047 7226 -537 7379
rect 4384 7324 4507 7379
rect 5453 16142 5460 16212
rect 5590 19689 12542 19716
rect 5590 19565 5662 19689
rect 12451 19565 12542 19689
rect 6985 19508 7113 19565
rect 10289 19508 10381 19565
rect 6985 19484 10381 19508
rect 5677 19339 6195 19374
rect 5677 19336 5907 19339
rect 5677 18103 5729 19336
rect 5891 19305 5907 19336
rect 6035 19305 6307 19339
rect 6435 19305 6707 19339
rect 6835 19305 7107 19339
rect 7235 19305 7507 19339
rect 7635 19305 7907 19339
rect 8035 19305 8307 19339
rect 8435 19305 8707 19339
rect 8835 19305 9107 19339
rect 9235 19305 9507 19339
rect 9635 19305 9907 19339
rect 10035 19305 10307 19339
rect 10435 19305 10707 19339
rect 10835 19305 11107 19339
rect 11235 19305 11507 19339
rect 11635 19305 11907 19339
rect 12035 19305 12051 19339
rect 5845 19255 5879 19271
rect 5845 18163 5879 18179
rect 6063 19255 6097 19271
rect 6063 18163 6097 18179
rect 6245 19255 6279 19271
rect 6245 18163 6279 18179
rect 6463 19255 6497 19271
rect 6463 18163 6497 18179
rect 6645 19255 6679 19271
rect 6645 18163 6679 18179
rect 6863 19255 6897 19271
rect 6863 18163 6897 18179
rect 7045 19255 7079 19271
rect 7045 18163 7079 18179
rect 7263 19255 7297 19271
rect 7263 18163 7297 18179
rect 7445 19255 7479 19271
rect 7445 18163 7479 18179
rect 7663 19255 7697 19271
rect 7663 18163 7697 18179
rect 7845 19255 7879 19271
rect 7845 18163 7879 18179
rect 8063 19255 8097 19271
rect 8063 18163 8097 18179
rect 8245 19255 8279 19271
rect 8245 18163 8279 18179
rect 8463 19255 8497 19271
rect 8463 18163 8497 18179
rect 8645 19255 8679 19271
rect 8645 18163 8679 18179
rect 8863 19255 8897 19271
rect 8863 18163 8897 18179
rect 9045 19255 9079 19271
rect 9045 18163 9079 18179
rect 9263 19255 9297 19271
rect 9263 18163 9297 18179
rect 9445 19255 9479 19271
rect 9445 18163 9479 18179
rect 9663 19255 9697 19271
rect 9663 18163 9697 18179
rect 9845 19255 9879 19271
rect 9845 18163 9879 18179
rect 10063 19255 10097 19271
rect 10063 18163 10097 18179
rect 10245 19255 10279 19271
rect 10245 18163 10279 18179
rect 10463 19255 10497 19271
rect 10463 18163 10497 18179
rect 10645 19255 10679 19271
rect 10645 18163 10679 18179
rect 10863 19255 10897 19271
rect 10863 18163 10897 18179
rect 11045 19255 11079 19271
rect 11045 18163 11079 18179
rect 11263 19255 11297 19271
rect 11263 18163 11297 18179
rect 11445 19255 11479 19271
rect 11445 18163 11479 18179
rect 11663 19255 11697 19271
rect 11663 18163 11697 18179
rect 11845 19255 11879 19271
rect 11845 18163 11879 18179
rect 12063 19255 12097 19271
rect 12063 18163 12097 18179
rect 5891 18103 5907 18129
rect 5677 18095 5907 18103
rect 6035 18095 6307 18129
rect 6435 18095 6707 18129
rect 6835 18095 7107 18129
rect 7235 18095 7507 18129
rect 7635 18095 7907 18129
rect 8035 18095 8307 18129
rect 8435 18095 8707 18129
rect 8835 18095 9107 18129
rect 9235 18095 9507 18129
rect 9635 18095 9907 18129
rect 10035 18095 10307 18129
rect 10435 18095 10707 18129
rect 10835 18095 11107 18129
rect 11235 18095 11507 18129
rect 11635 18095 11907 18129
rect 12035 18095 12051 18129
rect 5677 18065 6193 18095
rect 10074 17846 10247 18095
rect 10069 17815 10561 17846
rect 10069 17718 10110 17815
rect 10525 17718 10561 17815
rect 10069 17698 10561 17718
rect 8911 17676 8963 17677
rect 5770 17639 8963 17676
rect 5770 17605 5786 17639
rect 5914 17605 6186 17639
rect 6314 17605 6586 17639
rect 6714 17605 6986 17639
rect 7114 17605 7386 17639
rect 7514 17605 7786 17639
rect 7914 17605 8186 17639
rect 8314 17605 8586 17639
rect 8714 17628 8963 17639
rect 8714 17605 8730 17628
rect 5724 17555 5758 17571
rect 5724 16463 5758 16479
rect 5942 17555 5976 17571
rect 5942 16463 5976 16479
rect 6124 17555 6158 17571
rect 6124 16463 6158 16479
rect 6342 17555 6376 17571
rect 6342 16463 6376 16479
rect 6524 17555 6558 17571
rect 6524 16463 6558 16479
rect 6742 17555 6776 17571
rect 6742 16463 6776 16479
rect 6924 17555 6958 17571
rect 6924 16463 6958 16479
rect 7142 17555 7176 17571
rect 7142 16463 7176 16479
rect 7324 17555 7358 17571
rect 7324 16463 7358 16479
rect 7542 17555 7576 17571
rect 7542 16463 7576 16479
rect 7724 17555 7758 17571
rect 7724 16463 7758 16479
rect 7942 17555 7976 17571
rect 7942 16463 7976 16479
rect 8124 17555 8158 17571
rect 8124 16463 8158 16479
rect 8342 17555 8376 17571
rect 8342 16463 8376 16479
rect 8524 17555 8558 17571
rect 8524 16463 8558 16479
rect 8742 17555 8776 17571
rect 8742 16463 8776 16479
rect 5770 16395 5786 16429
rect 5914 16395 6186 16429
rect 6314 16395 6586 16429
rect 6714 16395 6986 16429
rect 7114 16395 7386 16429
rect 7514 16395 7786 16429
rect 7914 16395 8186 16429
rect 8314 16395 8586 16429
rect 8714 16410 8730 16429
rect 8911 16410 8963 17628
rect 9108 17585 9168 17619
rect 10222 17602 10282 17619
rect 10401 17602 10461 17608
rect 10222 17585 10461 17602
rect 9108 17559 9142 17585
rect 10248 17574 10461 17585
rect 12244 17574 12304 17608
rect 10248 17559 10435 17574
rect 9242 17418 9537 17419
rect 9229 17395 9537 17418
rect 9229 17377 9430 17395
rect 9229 17060 9274 17377
rect 9414 17361 9430 17377
rect 9558 17361 9830 17395
rect 9958 17361 9974 17395
rect 9368 17302 9402 17318
rect 9368 17110 9402 17126
rect 9586 17302 9620 17318
rect 9768 17302 9802 17318
rect 9620 17126 9768 17162
rect 9586 17112 9802 17126
rect 9586 17110 9620 17112
rect 9414 17060 9430 17067
rect 9229 17033 9430 17060
rect 9558 17033 9574 17067
rect 9229 17018 9551 17033
rect 9229 17016 9274 17018
rect 9108 16837 9142 16863
rect 9669 16837 9721 17112
rect 9768 17110 9802 17112
rect 9986 17302 10020 17318
rect 9986 17110 10020 17126
rect 9814 17033 9830 17067
rect 9958 17033 9974 17067
rect 10282 17548 10435 17559
rect 10282 16863 10401 17548
rect 10248 16837 10401 16863
rect 9108 16803 9168 16837
rect 10222 16824 10401 16837
rect 10222 16803 10282 16824
rect 12270 17548 12304 17574
rect 10673 17332 10689 17366
rect 10817 17332 11089 17366
rect 11217 17332 11489 17366
rect 11617 17332 11889 17366
rect 12017 17332 12033 17366
rect 10627 17273 10661 17289
rect 10627 17081 10661 17097
rect 10845 17273 10879 17289
rect 10845 17081 10879 17097
rect 10929 17038 10977 17332
rect 11027 17273 11061 17289
rect 11027 17081 11061 17097
rect 11245 17273 11279 17289
rect 11245 17081 11279 17097
rect 11427 17273 11461 17289
rect 11427 17081 11461 17097
rect 11645 17273 11679 17289
rect 11645 17081 11679 17097
rect 11725 17038 11773 17332
rect 11827 17273 11861 17289
rect 11827 17081 11861 17097
rect 12045 17273 12079 17289
rect 12045 17081 12079 17097
rect 10673 17004 10689 17038
rect 10817 17004 11089 17038
rect 11217 17004 11489 17038
rect 11617 17004 11889 17038
rect 12017 17004 12033 17038
rect 10401 16757 10435 16783
rect 11150 16851 11543 16867
rect 11150 16762 11180 16851
rect 11520 16762 11543 16851
rect 11150 16757 11543 16762
rect 12270 16757 12304 16783
rect 10401 16723 10461 16757
rect 12244 16723 12304 16757
rect 10509 16692 10811 16723
rect 9010 16473 9627 16505
rect 9010 16410 9052 16473
rect 8714 16395 9052 16410
rect 5770 16375 9052 16395
rect 9594 16375 9627 16473
rect 5770 16355 9627 16375
rect 9010 16343 9627 16355
rect 10509 16377 10546 16692
rect 10771 16377 10811 16692
rect 10509 16340 10811 16377
rect 6419 16266 8021 16293
rect 5590 16142 5655 16266
rect 12444 16142 12542 16266
rect 16247 18222 17282 19784
rect 5453 15720 8088 16142
rect 9336 15974 9683 16019
rect 8388 15720 8672 15725
rect 5453 15708 5734 15720
rect 4384 7226 4673 7324
rect 5452 15692 5734 15708
rect 5606 15630 5734 15692
rect 8648 15630 8672 15720
rect 9336 15686 9383 15974
rect 9629 15686 9683 15974
rect 10345 15720 10629 15725
rect 11510 15720 11938 16142
rect 12542 16126 12672 16142
rect 14352 18214 18330 18222
rect 14352 18198 14644 18214
rect 5606 15629 5849 15630
rect 8388 15625 8672 15630
rect 8861 15652 8921 15686
rect 10096 15652 10156 15686
rect 8861 15626 8895 15652
rect 5740 15521 7034 15557
rect 5740 15197 5782 15521
rect 5926 15487 5942 15521
rect 7018 15487 7034 15521
rect 7400 15477 8861 15523
rect 5858 15459 5892 15475
rect 5858 15315 5892 15331
rect 7068 15459 7102 15475
rect 7402 15443 7418 15477
rect 8494 15443 8510 15477
rect 7334 15415 7368 15431
rect 7334 15351 7368 15367
rect 8544 15415 8578 15431
rect 8544 15351 8578 15367
rect 7068 15315 7102 15331
rect 7238 15309 7278 15337
rect 7402 15309 7418 15339
rect 7238 15305 7418 15309
rect 8494 15305 8510 15339
rect 5926 15269 5942 15303
rect 7018 15269 7034 15303
rect 7238 15269 7622 15305
rect 5926 15233 7186 15269
rect 5740 15161 7034 15197
rect 5740 14837 5782 15161
rect 5926 15127 5942 15161
rect 7018 15127 7034 15161
rect 5858 15099 5892 15115
rect 5858 14955 5892 14971
rect 7068 15099 7102 15115
rect 7068 14955 7102 14971
rect 5926 14909 5942 14943
rect 7018 14909 7034 14943
rect 7150 14929 7186 15233
rect 7238 15015 7278 15269
rect 8640 15219 8680 15477
rect 7400 15179 8680 15219
rect 7400 15173 7418 15179
rect 7402 15145 7418 15173
rect 8494 15173 8680 15179
rect 8494 15145 8510 15173
rect 8730 15162 8802 15186
rect 7334 15117 7368 15133
rect 7334 15053 7368 15069
rect 8544 15117 8578 15133
rect 8544 15053 8578 15069
rect 8730 15079 8748 15162
rect 8783 15079 8802 15162
rect 7402 15015 7418 15041
rect 7238 15007 7418 15015
rect 8494 15007 8510 15041
rect 7238 14973 7670 15007
rect 8730 14948 8802 15079
rect 8298 14929 8802 14948
rect 7150 14912 8802 14929
rect 7150 14909 8480 14912
rect 5926 14897 8480 14909
rect 5926 14895 7388 14897
rect 5926 14873 7238 14895
rect 5740 14801 7034 14837
rect 5740 14477 5782 14801
rect 5926 14767 5942 14801
rect 7018 14767 7034 14801
rect 5858 14739 5892 14755
rect 5858 14595 5892 14611
rect 7068 14739 7102 14755
rect 7068 14595 7102 14611
rect 5926 14549 5942 14583
rect 7018 14549 7034 14583
rect 7178 14549 7238 14873
rect 7372 14863 7388 14895
rect 8464 14863 8480 14897
rect 7304 14835 7338 14851
rect 7304 14651 7338 14667
rect 8514 14835 8548 14851
rect 8514 14651 8548 14667
rect 7372 14605 7388 14639
rect 8464 14605 8480 14639
rect 7372 14571 8652 14605
rect 5926 14513 7238 14549
rect 7178 14507 7238 14513
rect 5740 14441 7034 14477
rect 5926 14407 5942 14441
rect 7018 14407 7034 14441
rect 7178 14473 8480 14507
rect 5858 14379 5892 14395
rect 5858 14235 5892 14251
rect 7068 14379 7102 14395
rect 7068 14235 7102 14251
rect 5926 14189 5942 14223
rect 7018 14189 7034 14223
rect 7178 14189 7220 14473
rect 7372 14439 7388 14473
rect 8464 14439 8480 14473
rect 7304 14411 7338 14427
rect 7304 14227 7338 14243
rect 8514 14411 8548 14427
rect 8514 14227 8548 14243
rect 8616 14305 8652 14571
rect 8616 14289 8759 14305
rect 5926 14153 7220 14189
rect 7372 14181 7388 14215
rect 8464 14185 8480 14215
rect 8616 14185 8641 14289
rect 8464 14181 8641 14185
rect 7372 14171 8641 14181
rect 7372 14156 8759 14171
rect 7442 14155 8759 14156
rect 7442 14151 8652 14155
rect 9336 15598 9383 15652
rect 9629 15598 9683 15652
rect 9336 15566 9433 15598
rect 9059 15518 9075 15552
rect 9251 15518 9267 15552
rect 8944 15490 9016 15506
rect 8944 15362 8982 15490
rect 8944 15346 9016 15362
rect 9310 15490 9381 15506
rect 9344 15362 9381 15490
rect 9310 15346 9381 15362
rect 8944 15220 8982 15346
rect 9059 15300 9075 15334
rect 9251 15300 9267 15334
rect 9344 15264 9381 15346
rect 9210 15242 9397 15264
rect 8944 15181 9115 15220
rect 9059 15144 9115 15181
rect 9210 15194 9274 15242
rect 9371 15194 9397 15242
rect 9210 15179 9397 15194
rect 9211 15144 9267 15179
rect 9059 15110 9075 15144
rect 9251 15110 9267 15144
rect 8982 15082 9016 15098
rect 8982 14828 9016 14954
rect 9310 15082 9344 15098
rect 9059 14892 9075 14926
rect 9251 14892 9267 14926
rect 9310 14851 9344 14954
rect 9271 14829 9376 14851
rect 9271 14828 9291 14829
rect 8982 14780 9291 14828
rect 8982 14636 9016 14780
rect 9271 14761 9291 14780
rect 9354 14761 9376 14829
rect 9271 14744 9376 14761
rect 9059 14664 9075 14698
rect 9251 14664 9267 14698
rect 8982 14252 9016 14268
rect 9310 14636 9344 14744
rect 9310 14252 9344 14268
rect 7442 14059 8428 14151
rect 8861 14126 8895 14152
rect 9058 14240 9268 14241
rect 9058 14206 9075 14240
rect 9251 14206 9268 14240
rect 9058 14126 9268 14206
rect 9467 14152 9550 15598
rect 9584 15566 9683 15598
rect 10122 15626 10156 15652
rect 9750 15518 9766 15552
rect 9942 15518 9958 15552
rect 9636 15490 9707 15506
rect 9636 15362 9673 15490
rect 9636 15346 9707 15362
rect 10001 15490 10073 15506
rect 10035 15362 10073 15490
rect 10001 15346 10073 15362
rect 9636 15264 9673 15346
rect 9750 15300 9766 15334
rect 9942 15300 9958 15334
rect 9620 15242 9807 15264
rect 9620 15194 9646 15242
rect 9743 15194 9807 15242
rect 10035 15220 10073 15346
rect 9620 15179 9807 15194
rect 9902 15181 10073 15220
rect 9750 15144 9806 15179
rect 9902 15144 9958 15181
rect 9750 15110 9766 15144
rect 9942 15110 9958 15144
rect 9673 15082 9707 15098
rect 9673 14851 9707 14954
rect 10001 15082 10035 15098
rect 9750 14892 9766 14926
rect 9942 14892 9958 14926
rect 9641 14829 9746 14851
rect 9641 14761 9663 14829
rect 9726 14828 9746 14829
rect 10001 14828 10035 14954
rect 9726 14780 10035 14828
rect 9726 14761 9746 14780
rect 9641 14744 9746 14761
rect 9673 14636 9707 14744
rect 9750 14664 9766 14698
rect 9942 14664 9958 14698
rect 9673 14252 9707 14268
rect 10001 14636 10035 14780
rect 10001 14252 10035 14268
rect 9433 14126 9584 14152
rect 9749 14240 9959 14241
rect 9749 14206 9766 14240
rect 9942 14206 9959 14240
rect 9749 14126 9959 14206
rect 10345 15630 10369 15720
rect 13283 15630 13299 15720
rect 13411 15692 13565 15708
rect 10345 15625 10629 15630
rect 10156 15477 11617 15523
rect 11983 15521 13277 15557
rect 11983 15487 11999 15521
rect 13075 15487 13091 15521
rect 10337 15219 10377 15477
rect 10507 15443 10523 15477
rect 11599 15443 11615 15477
rect 11915 15459 11949 15475
rect 10439 15415 10473 15431
rect 10439 15351 10473 15367
rect 11649 15415 11683 15431
rect 11649 15351 11683 15367
rect 10507 15305 10523 15339
rect 11599 15309 11615 15339
rect 11739 15309 11779 15337
rect 11915 15315 11949 15331
rect 13125 15459 13159 15475
rect 13125 15315 13159 15331
rect 11599 15305 11779 15309
rect 11395 15269 11779 15305
rect 11983 15269 11999 15303
rect 13075 15269 13091 15303
rect 10215 15162 10287 15186
rect 10337 15179 11617 15219
rect 10337 15173 10523 15179
rect 10215 15079 10234 15162
rect 10269 15079 10287 15162
rect 10507 15145 10523 15173
rect 11599 15173 11617 15179
rect 11599 15145 11615 15173
rect 10215 14948 10287 15079
rect 10439 15117 10473 15133
rect 10439 15053 10473 15069
rect 11649 15117 11683 15133
rect 11649 15053 11683 15069
rect 10507 15007 10523 15041
rect 11599 15015 11615 15041
rect 11739 15015 11779 15269
rect 11599 15007 11779 15015
rect 11347 14973 11779 15007
rect 11831 15233 13091 15269
rect 10215 14929 10719 14948
rect 11831 14929 11867 15233
rect 13235 15197 13277 15521
rect 11983 15161 13277 15197
rect 11983 15127 11999 15161
rect 13075 15127 13091 15161
rect 11915 15099 11949 15115
rect 11915 14955 11949 14971
rect 13125 15099 13159 15115
rect 13125 14955 13159 14971
rect 10215 14912 11867 14929
rect 10537 14909 11867 14912
rect 11983 14909 11999 14943
rect 13075 14909 13091 14943
rect 10537 14897 13091 14909
rect 10537 14863 10553 14897
rect 11629 14895 13091 14897
rect 11629 14863 11645 14895
rect 11779 14873 13091 14895
rect 10469 14835 10503 14851
rect 10469 14651 10503 14667
rect 11679 14835 11713 14851
rect 11679 14651 11713 14667
rect 10537 14605 10553 14639
rect 11629 14605 11645 14639
rect 10365 14571 11645 14605
rect 10365 14305 10401 14571
rect 11779 14549 11839 14873
rect 13235 14837 13277 15161
rect 11983 14801 13277 14837
rect 11983 14767 11999 14801
rect 13075 14767 13091 14801
rect 11915 14739 11949 14755
rect 11915 14595 11949 14611
rect 13125 14739 13159 14755
rect 13125 14595 13159 14611
rect 11983 14549 11999 14583
rect 13075 14549 13091 14583
rect 11779 14513 13091 14549
rect 11779 14507 11839 14513
rect 10537 14473 11839 14507
rect 13235 14477 13277 14801
rect 10537 14439 10553 14473
rect 11629 14439 11645 14473
rect 10258 14289 10401 14305
rect 10376 14185 10401 14289
rect 10469 14411 10503 14427
rect 10469 14227 10503 14243
rect 11679 14411 11713 14427
rect 11679 14227 11713 14243
rect 10537 14185 10553 14215
rect 10376 14181 10553 14185
rect 11629 14181 11645 14215
rect 10376 14171 11645 14181
rect 10258 14156 11645 14171
rect 11797 14189 11839 14473
rect 11983 14441 13277 14477
rect 11983 14407 11999 14441
rect 13075 14407 13091 14441
rect 11915 14379 11949 14395
rect 11915 14235 11949 14251
rect 13125 14379 13159 14395
rect 13125 14235 13159 14251
rect 11983 14189 11999 14223
rect 13075 14189 13091 14223
rect 10258 14155 11575 14156
rect 10122 14126 10156 14152
rect 10365 14151 11575 14155
rect 11797 14153 13091 14189
rect 8861 14092 8921 14126
rect 9407 14092 9610 14126
rect 10096 14092 10156 14126
rect 7442 14054 8672 14059
rect 5718 13964 5734 14054
rect 8648 13964 8672 14054
rect 9467 14020 9550 14092
rect 10589 14059 11575 14151
rect 10345 14054 11575 14059
rect 8388 13959 8672 13964
rect 8861 13986 8921 14020
rect 9407 13986 9610 14020
rect 10096 13986 10156 14020
rect 8861 13960 8895 13986
rect 5740 13855 7034 13891
rect 5740 13531 5782 13855
rect 5926 13821 5942 13855
rect 7018 13821 7034 13855
rect 7400 13811 8861 13857
rect 5858 13793 5892 13809
rect 5858 13649 5892 13665
rect 7068 13793 7102 13809
rect 7402 13777 7418 13811
rect 8494 13777 8510 13811
rect 7334 13749 7368 13765
rect 7334 13685 7368 13701
rect 8544 13749 8578 13765
rect 8544 13685 8578 13701
rect 7068 13649 7102 13665
rect 7238 13643 7278 13671
rect 7402 13643 7418 13673
rect 7238 13639 7418 13643
rect 8494 13639 8510 13673
rect 5926 13603 5942 13637
rect 7018 13603 7034 13637
rect 7238 13603 7622 13639
rect 5926 13567 7186 13603
rect 5740 13495 7034 13531
rect 5740 13171 5782 13495
rect 5926 13461 5942 13495
rect 7018 13461 7034 13495
rect 5858 13433 5892 13449
rect 5858 13289 5892 13305
rect 7068 13433 7102 13449
rect 7068 13289 7102 13305
rect 5926 13243 5942 13277
rect 7018 13243 7034 13277
rect 7150 13263 7186 13567
rect 7238 13349 7278 13603
rect 8640 13553 8680 13811
rect 7400 13513 8680 13553
rect 7400 13507 7418 13513
rect 7402 13479 7418 13507
rect 8494 13507 8680 13513
rect 8494 13479 8510 13507
rect 8730 13496 8802 13520
rect 7334 13451 7368 13467
rect 7334 13387 7368 13403
rect 8544 13451 8578 13467
rect 8544 13387 8578 13403
rect 8730 13413 8748 13496
rect 8783 13413 8802 13496
rect 7402 13349 7418 13375
rect 7238 13341 7418 13349
rect 8494 13341 8510 13375
rect 7238 13307 7670 13341
rect 8730 13282 8802 13413
rect 8298 13263 8802 13282
rect 7150 13246 8802 13263
rect 7150 13243 8480 13246
rect 5926 13231 8480 13243
rect 5926 13229 7388 13231
rect 5926 13207 7238 13229
rect 5740 13135 7034 13171
rect 5740 12811 5782 13135
rect 5926 13101 5942 13135
rect 7018 13101 7034 13135
rect 5858 13073 5892 13089
rect 5858 12929 5892 12945
rect 7068 13073 7102 13089
rect 7068 12929 7102 12945
rect 5926 12883 5942 12917
rect 7018 12883 7034 12917
rect 7178 12883 7238 13207
rect 7372 13197 7388 13229
rect 8464 13197 8480 13231
rect 7304 13169 7338 13185
rect 7304 12985 7338 13001
rect 8514 13169 8548 13185
rect 8514 12985 8548 13001
rect 7372 12939 7388 12973
rect 8464 12939 8480 12973
rect 7372 12905 8652 12939
rect 5926 12847 7238 12883
rect 7178 12841 7238 12847
rect 5740 12775 7034 12811
rect 5926 12741 5942 12775
rect 7018 12741 7034 12775
rect 7178 12807 8480 12841
rect 5858 12713 5892 12729
rect 5858 12569 5892 12585
rect 7068 12713 7102 12729
rect 7068 12569 7102 12585
rect 5926 12523 5942 12557
rect 7018 12523 7034 12557
rect 7178 12523 7220 12807
rect 7372 12773 7388 12807
rect 8464 12773 8480 12807
rect 7304 12745 7338 12761
rect 7304 12561 7338 12577
rect 8514 12745 8548 12761
rect 8514 12561 8548 12577
rect 8616 12639 8652 12905
rect 8616 12623 8759 12639
rect 5926 12487 7220 12523
rect 7372 12515 7388 12549
rect 8464 12519 8480 12549
rect 8616 12519 8641 12623
rect 8464 12515 8641 12519
rect 7372 12505 8641 12515
rect 7372 12490 8759 12505
rect 7442 12489 8759 12490
rect 7442 12485 8652 12489
rect 9336 13960 9681 13986
rect 9336 13902 9433 13960
rect 9059 13852 9075 13886
rect 9251 13852 9267 13886
rect 8944 13824 9016 13840
rect 8944 13696 8982 13824
rect 8944 13680 9016 13696
rect 9310 13824 9381 13840
rect 9344 13696 9381 13824
rect 9310 13680 9381 13696
rect 8944 13554 8982 13680
rect 9059 13634 9075 13668
rect 9251 13634 9267 13668
rect 9344 13598 9381 13680
rect 9210 13576 9397 13598
rect 8944 13515 9115 13554
rect 9059 13478 9115 13515
rect 9210 13528 9274 13576
rect 9371 13528 9397 13576
rect 9210 13513 9397 13528
rect 9211 13478 9267 13513
rect 9059 13444 9075 13478
rect 9251 13444 9267 13478
rect 8982 13416 9016 13432
rect 8982 13162 9016 13288
rect 9310 13416 9344 13432
rect 9059 13226 9075 13260
rect 9251 13226 9267 13260
rect 9310 13185 9344 13288
rect 9271 13163 9376 13185
rect 9271 13162 9291 13163
rect 8982 13114 9291 13162
rect 8982 12970 9016 13114
rect 9271 13095 9291 13114
rect 9354 13095 9376 13163
rect 9271 13078 9376 13095
rect 9059 12998 9075 13032
rect 9251 12998 9267 13032
rect 8982 12586 9016 12602
rect 9310 12970 9344 13078
rect 9310 12586 9344 12602
rect 7442 12393 8428 12485
rect 8861 12460 8895 12486
rect 9058 12574 9268 12575
rect 9058 12540 9075 12574
rect 9251 12540 9268 12574
rect 9058 12460 9268 12540
rect 9467 12486 9550 13960
rect 9584 13902 9681 13960
rect 10122 13960 10156 13986
rect 9750 13852 9766 13886
rect 9942 13852 9958 13886
rect 9636 13824 9707 13840
rect 9636 13696 9673 13824
rect 9636 13680 9707 13696
rect 10001 13824 10073 13840
rect 10035 13696 10073 13824
rect 10001 13680 10073 13696
rect 9636 13598 9673 13680
rect 9750 13634 9766 13668
rect 9942 13634 9958 13668
rect 9620 13576 9807 13598
rect 9620 13528 9646 13576
rect 9743 13528 9807 13576
rect 10035 13554 10073 13680
rect 9620 13513 9807 13528
rect 9902 13515 10073 13554
rect 9750 13478 9806 13513
rect 9902 13478 9958 13515
rect 9750 13444 9766 13478
rect 9942 13444 9958 13478
rect 9673 13416 9707 13432
rect 9673 13185 9707 13288
rect 10001 13416 10035 13432
rect 9750 13226 9766 13260
rect 9942 13226 9958 13260
rect 9641 13163 9746 13185
rect 9641 13095 9663 13163
rect 9726 13162 9746 13163
rect 10001 13162 10035 13288
rect 9726 13114 10035 13162
rect 9726 13095 9746 13114
rect 9641 13078 9746 13095
rect 9673 12970 9707 13078
rect 9750 12998 9766 13032
rect 9942 12998 9958 13032
rect 9673 12586 9707 12602
rect 10001 12970 10035 13114
rect 10001 12586 10035 12602
rect 9433 12460 9584 12486
rect 9749 12574 9959 12575
rect 9749 12540 9766 12574
rect 9942 12540 9959 12574
rect 9749 12460 9959 12540
rect 10345 13964 10369 14054
rect 13283 13964 13299 14054
rect 10345 13959 10629 13964
rect 10156 13811 11617 13857
rect 11983 13855 13277 13891
rect 11983 13821 11999 13855
rect 13075 13821 13091 13855
rect 10337 13553 10377 13811
rect 10507 13777 10523 13811
rect 11599 13777 11615 13811
rect 11915 13793 11949 13809
rect 10439 13749 10473 13765
rect 10439 13685 10473 13701
rect 11649 13749 11683 13765
rect 11649 13685 11683 13701
rect 10507 13639 10523 13673
rect 11599 13643 11615 13673
rect 11739 13643 11779 13671
rect 11915 13649 11949 13665
rect 13125 13793 13159 13809
rect 13125 13649 13159 13665
rect 11599 13639 11779 13643
rect 11395 13603 11779 13639
rect 11983 13603 11999 13637
rect 13075 13603 13091 13637
rect 10215 13496 10287 13520
rect 10337 13513 11617 13553
rect 10337 13507 10523 13513
rect 10215 13413 10234 13496
rect 10269 13413 10287 13496
rect 10507 13479 10523 13507
rect 11599 13507 11617 13513
rect 11599 13479 11615 13507
rect 10215 13282 10287 13413
rect 10439 13451 10473 13467
rect 10439 13387 10473 13403
rect 11649 13451 11683 13467
rect 11649 13387 11683 13403
rect 10507 13341 10523 13375
rect 11599 13349 11615 13375
rect 11739 13349 11779 13603
rect 11599 13341 11779 13349
rect 11347 13307 11779 13341
rect 11831 13567 13091 13603
rect 10215 13263 10719 13282
rect 11831 13263 11867 13567
rect 13235 13531 13277 13855
rect 11983 13495 13277 13531
rect 11983 13461 11999 13495
rect 13075 13461 13091 13495
rect 11915 13433 11949 13449
rect 11915 13289 11949 13305
rect 13125 13433 13159 13449
rect 13125 13289 13159 13305
rect 10215 13246 11867 13263
rect 10537 13243 11867 13246
rect 11983 13243 11999 13277
rect 13075 13243 13091 13277
rect 10537 13231 13091 13243
rect 10537 13197 10553 13231
rect 11629 13229 13091 13231
rect 11629 13197 11645 13229
rect 11779 13207 13091 13229
rect 10469 13169 10503 13185
rect 10469 12985 10503 13001
rect 11679 13169 11713 13185
rect 11679 12985 11713 13001
rect 10537 12939 10553 12973
rect 11629 12939 11645 12973
rect 10365 12905 11645 12939
rect 10365 12639 10401 12905
rect 11779 12883 11839 13207
rect 13235 13171 13277 13495
rect 11983 13135 13277 13171
rect 11983 13101 11999 13135
rect 13075 13101 13091 13135
rect 11915 13073 11949 13089
rect 11915 12929 11949 12945
rect 13125 13073 13159 13089
rect 13125 12929 13159 12945
rect 11983 12883 11999 12917
rect 13075 12883 13091 12917
rect 11779 12847 13091 12883
rect 11779 12841 11839 12847
rect 10537 12807 11839 12841
rect 13235 12811 13277 13135
rect 10537 12773 10553 12807
rect 11629 12773 11645 12807
rect 10258 12623 10401 12639
rect 10376 12519 10401 12623
rect 10469 12745 10503 12761
rect 10469 12561 10503 12577
rect 11679 12745 11713 12761
rect 11679 12561 11713 12577
rect 10537 12519 10553 12549
rect 10376 12515 10553 12519
rect 11629 12515 11645 12549
rect 10376 12505 11645 12515
rect 10258 12490 11645 12505
rect 11797 12523 11839 12807
rect 11983 12775 13277 12811
rect 11983 12741 11999 12775
rect 13075 12741 13091 12775
rect 11915 12713 11949 12729
rect 11915 12569 11949 12585
rect 13125 12713 13159 12729
rect 13125 12569 13159 12585
rect 11983 12523 11999 12557
rect 13075 12523 13091 12557
rect 10258 12489 11575 12490
rect 10122 12460 10156 12486
rect 10365 12485 11575 12489
rect 11797 12487 13091 12523
rect 8861 12426 8921 12460
rect 9407 12426 9610 12460
rect 10096 12426 10156 12460
rect 7442 12388 8672 12393
rect 5718 12298 5734 12388
rect 8648 12298 8672 12388
rect 9467 12354 9550 12426
rect 10589 12393 11575 12485
rect 10345 12388 11575 12393
rect 8388 12293 8672 12298
rect 8861 12320 8921 12354
rect 9407 12320 9610 12354
rect 10096 12320 10156 12354
rect 8861 12294 8895 12320
rect 5740 12189 7034 12225
rect 5740 11865 5782 12189
rect 5926 12155 5942 12189
rect 7018 12155 7034 12189
rect 7400 12145 8861 12191
rect 5858 12127 5892 12143
rect 5858 11983 5892 11999
rect 7068 12127 7102 12143
rect 7402 12111 7418 12145
rect 8494 12111 8510 12145
rect 7334 12083 7368 12099
rect 7334 12019 7368 12035
rect 8544 12083 8578 12099
rect 8544 12019 8578 12035
rect 7068 11983 7102 11999
rect 7238 11977 7278 12005
rect 7402 11977 7418 12007
rect 7238 11973 7418 11977
rect 8494 11973 8510 12007
rect 5926 11937 5942 11971
rect 7018 11937 7034 11971
rect 7238 11937 7622 11973
rect 5926 11901 7186 11937
rect 5740 11829 7034 11865
rect 5740 11505 5782 11829
rect 5926 11795 5942 11829
rect 7018 11795 7034 11829
rect 5858 11767 5892 11783
rect 5858 11623 5892 11639
rect 7068 11767 7102 11783
rect 7068 11623 7102 11639
rect 5926 11577 5942 11611
rect 7018 11577 7034 11611
rect 7150 11597 7186 11901
rect 7238 11683 7278 11937
rect 8640 11887 8680 12145
rect 7400 11847 8680 11887
rect 7400 11841 7418 11847
rect 7402 11813 7418 11841
rect 8494 11841 8680 11847
rect 8494 11813 8510 11841
rect 8730 11830 8802 11854
rect 7334 11785 7368 11801
rect 7334 11721 7368 11737
rect 8544 11785 8578 11801
rect 8544 11721 8578 11737
rect 8730 11747 8748 11830
rect 8783 11747 8802 11830
rect 7402 11683 7418 11709
rect 7238 11675 7418 11683
rect 8494 11675 8510 11709
rect 7238 11641 7670 11675
rect 8730 11616 8802 11747
rect 8298 11597 8802 11616
rect 7150 11580 8802 11597
rect 7150 11577 8480 11580
rect 5926 11565 8480 11577
rect 5926 11563 7388 11565
rect 5926 11541 7238 11563
rect 5740 11469 7034 11505
rect 5740 11145 5782 11469
rect 5926 11435 5942 11469
rect 7018 11435 7034 11469
rect 5858 11407 5892 11423
rect 5858 11263 5892 11279
rect 7068 11407 7102 11423
rect 7068 11263 7102 11279
rect 5926 11217 5942 11251
rect 7018 11217 7034 11251
rect 7178 11217 7238 11541
rect 7372 11531 7388 11563
rect 8464 11531 8480 11565
rect 7304 11503 7338 11519
rect 7304 11319 7338 11335
rect 8514 11503 8548 11519
rect 8514 11319 8548 11335
rect 7372 11273 7388 11307
rect 8464 11273 8480 11307
rect 7372 11239 8652 11273
rect 5926 11181 7238 11217
rect 7178 11175 7238 11181
rect 5740 11109 7034 11145
rect 5926 11075 5942 11109
rect 7018 11075 7034 11109
rect 7178 11141 8480 11175
rect 5858 11047 5892 11063
rect 5858 10903 5892 10919
rect 7068 11047 7102 11063
rect 7068 10903 7102 10919
rect 5926 10857 5942 10891
rect 7018 10857 7034 10891
rect 7178 10857 7220 11141
rect 7372 11107 7388 11141
rect 8464 11107 8480 11141
rect 7304 11079 7338 11095
rect 7304 10895 7338 10911
rect 8514 11079 8548 11095
rect 8514 10895 8548 10911
rect 8616 10973 8652 11239
rect 8616 10957 8759 10973
rect 5926 10821 7220 10857
rect 7372 10849 7388 10883
rect 8464 10853 8480 10883
rect 8616 10853 8641 10957
rect 8464 10849 8641 10853
rect 7372 10839 8641 10849
rect 7372 10824 8759 10839
rect 7442 10823 8759 10824
rect 7442 10819 8652 10823
rect 9336 12294 9681 12320
rect 9336 12236 9433 12294
rect 9059 12186 9075 12220
rect 9251 12186 9267 12220
rect 8944 12158 9016 12174
rect 8944 12030 8982 12158
rect 8944 12014 9016 12030
rect 9310 12158 9381 12174
rect 9344 12030 9381 12158
rect 9310 12014 9381 12030
rect 8944 11888 8982 12014
rect 9059 11968 9075 12002
rect 9251 11968 9267 12002
rect 9344 11932 9381 12014
rect 9210 11910 9397 11932
rect 8944 11849 9115 11888
rect 9059 11812 9115 11849
rect 9210 11862 9274 11910
rect 9371 11862 9397 11910
rect 9210 11847 9397 11862
rect 9211 11812 9267 11847
rect 9059 11778 9075 11812
rect 9251 11778 9267 11812
rect 8982 11750 9016 11766
rect 8982 11496 9016 11622
rect 9310 11750 9344 11766
rect 9059 11560 9075 11594
rect 9251 11560 9267 11594
rect 9310 11519 9344 11622
rect 9271 11497 9376 11519
rect 9271 11496 9291 11497
rect 8982 11448 9291 11496
rect 8982 11304 9016 11448
rect 9271 11429 9291 11448
rect 9354 11429 9376 11497
rect 9271 11412 9376 11429
rect 9059 11332 9075 11366
rect 9251 11332 9267 11366
rect 8982 10920 9016 10936
rect 9310 11304 9344 11412
rect 9310 10920 9344 10936
rect 7442 10727 8428 10819
rect 8861 10794 8895 10820
rect 9058 10908 9268 10909
rect 9058 10874 9075 10908
rect 9251 10874 9268 10908
rect 9058 10794 9268 10874
rect 9467 10820 9550 12294
rect 9584 12236 9681 12294
rect 10122 12294 10156 12320
rect 9750 12186 9766 12220
rect 9942 12186 9958 12220
rect 9636 12158 9707 12174
rect 9636 12030 9673 12158
rect 9636 12014 9707 12030
rect 10001 12158 10073 12174
rect 10035 12030 10073 12158
rect 10001 12014 10073 12030
rect 9636 11932 9673 12014
rect 9750 11968 9766 12002
rect 9942 11968 9958 12002
rect 9620 11910 9807 11932
rect 9620 11862 9646 11910
rect 9743 11862 9807 11910
rect 10035 11888 10073 12014
rect 9620 11847 9807 11862
rect 9902 11849 10073 11888
rect 9750 11812 9806 11847
rect 9902 11812 9958 11849
rect 9750 11778 9766 11812
rect 9942 11778 9958 11812
rect 9673 11750 9707 11766
rect 9673 11519 9707 11622
rect 10001 11750 10035 11766
rect 9750 11560 9766 11594
rect 9942 11560 9958 11594
rect 9641 11497 9746 11519
rect 9641 11429 9663 11497
rect 9726 11496 9746 11497
rect 10001 11496 10035 11622
rect 9726 11448 10035 11496
rect 9726 11429 9746 11448
rect 9641 11412 9746 11429
rect 9673 11304 9707 11412
rect 9750 11332 9766 11366
rect 9942 11332 9958 11366
rect 9673 10920 9707 10936
rect 10001 11304 10035 11448
rect 10001 10920 10035 10936
rect 9433 10794 9584 10820
rect 9749 10908 9959 10909
rect 9749 10874 9766 10908
rect 9942 10874 9959 10908
rect 9749 10794 9959 10874
rect 10345 12298 10369 12388
rect 13283 12298 13299 12388
rect 10345 12293 10629 12298
rect 10156 12145 11617 12191
rect 11983 12189 13277 12225
rect 11983 12155 11999 12189
rect 13075 12155 13091 12189
rect 10337 11887 10377 12145
rect 10507 12111 10523 12145
rect 11599 12111 11615 12145
rect 11915 12127 11949 12143
rect 10439 12083 10473 12099
rect 10439 12019 10473 12035
rect 11649 12083 11683 12099
rect 11649 12019 11683 12035
rect 10507 11973 10523 12007
rect 11599 11977 11615 12007
rect 11739 11977 11779 12005
rect 11915 11983 11949 11999
rect 13125 12127 13159 12143
rect 13125 11983 13159 11999
rect 11599 11973 11779 11977
rect 11395 11937 11779 11973
rect 11983 11937 11999 11971
rect 13075 11937 13091 11971
rect 10215 11830 10287 11854
rect 10337 11847 11617 11887
rect 10337 11841 10523 11847
rect 10215 11747 10234 11830
rect 10269 11747 10287 11830
rect 10507 11813 10523 11841
rect 11599 11841 11617 11847
rect 11599 11813 11615 11841
rect 10215 11616 10287 11747
rect 10439 11785 10473 11801
rect 10439 11721 10473 11737
rect 11649 11785 11683 11801
rect 11649 11721 11683 11737
rect 10507 11675 10523 11709
rect 11599 11683 11615 11709
rect 11739 11683 11779 11937
rect 11599 11675 11779 11683
rect 11347 11641 11779 11675
rect 11831 11901 13091 11937
rect 10215 11597 10719 11616
rect 11831 11597 11867 11901
rect 13235 11865 13277 12189
rect 11983 11829 13277 11865
rect 11983 11795 11999 11829
rect 13075 11795 13091 11829
rect 11915 11767 11949 11783
rect 11915 11623 11949 11639
rect 13125 11767 13159 11783
rect 13125 11623 13159 11639
rect 10215 11580 11867 11597
rect 10537 11577 11867 11580
rect 11983 11577 11999 11611
rect 13075 11577 13091 11611
rect 10537 11565 13091 11577
rect 10537 11531 10553 11565
rect 11629 11563 13091 11565
rect 11629 11531 11645 11563
rect 11779 11541 13091 11563
rect 10469 11503 10503 11519
rect 10469 11319 10503 11335
rect 11679 11503 11713 11519
rect 11679 11319 11713 11335
rect 10537 11273 10553 11307
rect 11629 11273 11645 11307
rect 10365 11239 11645 11273
rect 10365 10973 10401 11239
rect 11779 11217 11839 11541
rect 13235 11505 13277 11829
rect 11983 11469 13277 11505
rect 11983 11435 11999 11469
rect 13075 11435 13091 11469
rect 11915 11407 11949 11423
rect 11915 11263 11949 11279
rect 13125 11407 13159 11423
rect 13125 11263 13159 11279
rect 11983 11217 11999 11251
rect 13075 11217 13091 11251
rect 11779 11181 13091 11217
rect 11779 11175 11839 11181
rect 10537 11141 11839 11175
rect 13235 11145 13277 11469
rect 10537 11107 10553 11141
rect 11629 11107 11645 11141
rect 10258 10957 10401 10973
rect 10376 10853 10401 10957
rect 10469 11079 10503 11095
rect 10469 10895 10503 10911
rect 11679 11079 11713 11095
rect 11679 10895 11713 10911
rect 10537 10853 10553 10883
rect 10376 10849 10553 10853
rect 11629 10849 11645 10883
rect 10376 10839 11645 10849
rect 10258 10824 11645 10839
rect 11797 10857 11839 11141
rect 11983 11109 13277 11145
rect 11983 11075 11999 11109
rect 13075 11075 13091 11109
rect 11915 11047 11949 11063
rect 11915 10903 11949 10919
rect 13125 11047 13159 11063
rect 13125 10903 13159 10919
rect 11983 10857 11999 10891
rect 13075 10857 13091 10891
rect 10258 10823 11575 10824
rect 10122 10794 10156 10820
rect 10365 10819 11575 10823
rect 11797 10821 13091 10857
rect 8861 10760 8921 10794
rect 9407 10760 9610 10794
rect 10096 10760 10156 10794
rect 7442 10722 8672 10727
rect 5718 10632 5734 10722
rect 8648 10632 8672 10722
rect 9467 10688 9550 10760
rect 10589 10727 11575 10819
rect 10345 10722 11575 10727
rect 8388 10627 8672 10632
rect 8861 10654 8921 10688
rect 9407 10654 9610 10688
rect 10096 10654 10156 10688
rect 8861 10628 8895 10654
rect 5740 10523 7034 10559
rect 5740 10199 5782 10523
rect 5926 10489 5942 10523
rect 7018 10489 7034 10523
rect 7400 10479 8861 10525
rect 5858 10461 5892 10477
rect 5858 10317 5892 10333
rect 7068 10461 7102 10477
rect 7402 10445 7418 10479
rect 8494 10445 8510 10479
rect 7334 10417 7368 10433
rect 7334 10353 7368 10369
rect 8544 10417 8578 10433
rect 8544 10353 8578 10369
rect 7068 10317 7102 10333
rect 7238 10311 7278 10339
rect 7402 10311 7418 10341
rect 7238 10307 7418 10311
rect 8494 10307 8510 10341
rect 5926 10271 5942 10305
rect 7018 10271 7034 10305
rect 7238 10271 7622 10307
rect 5926 10235 7186 10271
rect 5740 10163 7034 10199
rect 5740 9839 5782 10163
rect 5926 10129 5942 10163
rect 7018 10129 7034 10163
rect 5858 10101 5892 10117
rect 5858 9957 5892 9973
rect 7068 10101 7102 10117
rect 7068 9957 7102 9973
rect 5926 9911 5942 9945
rect 7018 9911 7034 9945
rect 7150 9931 7186 10235
rect 7238 10017 7278 10271
rect 8640 10221 8680 10479
rect 7400 10181 8680 10221
rect 7400 10175 7418 10181
rect 7402 10147 7418 10175
rect 8494 10175 8680 10181
rect 8494 10147 8510 10175
rect 8730 10164 8802 10188
rect 7334 10119 7368 10135
rect 7334 10055 7368 10071
rect 8544 10119 8578 10135
rect 8544 10055 8578 10071
rect 8730 10081 8748 10164
rect 8783 10081 8802 10164
rect 7402 10017 7418 10043
rect 7238 10009 7418 10017
rect 8494 10009 8510 10043
rect 7238 9975 7670 10009
rect 8730 9950 8802 10081
rect 8298 9931 8802 9950
rect 7150 9914 8802 9931
rect 7150 9911 8480 9914
rect 5926 9899 8480 9911
rect 5926 9897 7388 9899
rect 5926 9875 7238 9897
rect 5740 9803 7034 9839
rect 5740 9479 5782 9803
rect 5926 9769 5942 9803
rect 7018 9769 7034 9803
rect 5858 9741 5892 9757
rect 5858 9597 5892 9613
rect 7068 9741 7102 9757
rect 7068 9597 7102 9613
rect 5926 9551 5942 9585
rect 7018 9551 7034 9585
rect 7178 9551 7238 9875
rect 7372 9865 7388 9897
rect 8464 9865 8480 9899
rect 7304 9837 7338 9853
rect 7304 9653 7338 9669
rect 8514 9837 8548 9853
rect 8514 9653 8548 9669
rect 7372 9607 7388 9641
rect 8464 9607 8480 9641
rect 7372 9573 8652 9607
rect 5926 9515 7238 9551
rect 7178 9509 7238 9515
rect 5740 9443 7034 9479
rect 5926 9409 5942 9443
rect 7018 9409 7034 9443
rect 7178 9475 8480 9509
rect 5858 9381 5892 9397
rect 5858 9237 5892 9253
rect 7068 9381 7102 9397
rect 7068 9237 7102 9253
rect 5926 9191 5942 9225
rect 7018 9191 7034 9225
rect 7178 9191 7220 9475
rect 7372 9441 7388 9475
rect 8464 9441 8480 9475
rect 7304 9413 7338 9429
rect 7304 9229 7338 9245
rect 8514 9413 8548 9429
rect 8514 9229 8548 9245
rect 8616 9307 8652 9573
rect 8616 9291 8759 9307
rect 5926 9155 7220 9191
rect 7372 9183 7388 9217
rect 8464 9187 8480 9217
rect 8616 9187 8641 9291
rect 8464 9183 8641 9187
rect 7372 9173 8641 9183
rect 7372 9158 8759 9173
rect 7442 9157 8759 9158
rect 7442 9153 8652 9157
rect 9336 10628 9681 10654
rect 9336 10570 9433 10628
rect 9059 10520 9075 10554
rect 9251 10520 9267 10554
rect 8944 10492 9016 10508
rect 8944 10364 8982 10492
rect 8944 10348 9016 10364
rect 9310 10492 9381 10508
rect 9344 10364 9381 10492
rect 9310 10348 9381 10364
rect 8944 10222 8982 10348
rect 9059 10302 9075 10336
rect 9251 10302 9267 10336
rect 9344 10266 9381 10348
rect 9210 10244 9397 10266
rect 8944 10183 9115 10222
rect 9059 10146 9115 10183
rect 9210 10196 9274 10244
rect 9371 10196 9397 10244
rect 9210 10181 9397 10196
rect 9211 10146 9267 10181
rect 9059 10112 9075 10146
rect 9251 10112 9267 10146
rect 8982 10084 9016 10100
rect 8982 9830 9016 9956
rect 9310 10084 9344 10100
rect 9059 9894 9075 9928
rect 9251 9894 9267 9928
rect 9310 9853 9344 9956
rect 9271 9831 9376 9853
rect 9271 9830 9291 9831
rect 8982 9782 9291 9830
rect 8982 9638 9016 9782
rect 9271 9763 9291 9782
rect 9354 9763 9376 9831
rect 9271 9746 9376 9763
rect 9059 9666 9075 9700
rect 9251 9666 9267 9700
rect 8982 9254 9016 9270
rect 9310 9638 9344 9746
rect 9310 9254 9344 9270
rect 7442 9061 8428 9153
rect 8861 9128 8895 9154
rect 9058 9242 9268 9243
rect 9058 9208 9075 9242
rect 9251 9208 9268 9242
rect 9058 9128 9268 9208
rect 9467 9154 9550 10628
rect 9584 10570 9681 10628
rect 10122 10628 10156 10654
rect 9750 10520 9766 10554
rect 9942 10520 9958 10554
rect 9636 10492 9707 10508
rect 9636 10364 9673 10492
rect 9636 10348 9707 10364
rect 10001 10492 10073 10508
rect 10035 10364 10073 10492
rect 10001 10348 10073 10364
rect 9636 10266 9673 10348
rect 9750 10302 9766 10336
rect 9942 10302 9958 10336
rect 9620 10244 9807 10266
rect 9620 10196 9646 10244
rect 9743 10196 9807 10244
rect 10035 10222 10073 10348
rect 9620 10181 9807 10196
rect 9902 10183 10073 10222
rect 9750 10146 9806 10181
rect 9902 10146 9958 10183
rect 9750 10112 9766 10146
rect 9942 10112 9958 10146
rect 9673 10084 9707 10100
rect 9673 9853 9707 9956
rect 10001 10084 10035 10100
rect 9750 9894 9766 9928
rect 9942 9894 9958 9928
rect 9641 9831 9746 9853
rect 9641 9763 9663 9831
rect 9726 9830 9746 9831
rect 10001 9830 10035 9956
rect 9726 9782 10035 9830
rect 9726 9763 9746 9782
rect 9641 9746 9746 9763
rect 9673 9638 9707 9746
rect 9750 9666 9766 9700
rect 9942 9666 9958 9700
rect 9673 9254 9707 9270
rect 10001 9638 10035 9782
rect 10001 9254 10035 9270
rect 9433 9128 9584 9154
rect 9749 9242 9959 9243
rect 9749 9208 9766 9242
rect 9942 9208 9959 9242
rect 9749 9128 9959 9208
rect 10345 10632 10369 10722
rect 13283 10632 13299 10722
rect 10345 10627 10629 10632
rect 10156 10479 11617 10525
rect 11983 10523 13277 10559
rect 11983 10489 11999 10523
rect 13075 10489 13091 10523
rect 10337 10221 10377 10479
rect 10507 10445 10523 10479
rect 11599 10445 11615 10479
rect 11915 10461 11949 10477
rect 10439 10417 10473 10433
rect 10439 10353 10473 10369
rect 11649 10417 11683 10433
rect 11649 10353 11683 10369
rect 10507 10307 10523 10341
rect 11599 10311 11615 10341
rect 11739 10311 11779 10339
rect 11915 10317 11949 10333
rect 13125 10461 13159 10477
rect 13125 10317 13159 10333
rect 11599 10307 11779 10311
rect 11395 10271 11779 10307
rect 11983 10271 11999 10305
rect 13075 10271 13091 10305
rect 10215 10164 10287 10188
rect 10337 10181 11617 10221
rect 10337 10175 10523 10181
rect 10215 10081 10234 10164
rect 10269 10081 10287 10164
rect 10507 10147 10523 10175
rect 11599 10175 11617 10181
rect 11599 10147 11615 10175
rect 10215 9950 10287 10081
rect 10439 10119 10473 10135
rect 10439 10055 10473 10071
rect 11649 10119 11683 10135
rect 11649 10055 11683 10071
rect 10507 10009 10523 10043
rect 11599 10017 11615 10043
rect 11739 10017 11779 10271
rect 11599 10009 11779 10017
rect 11347 9975 11779 10009
rect 11831 10235 13091 10271
rect 10215 9931 10719 9950
rect 11831 9931 11867 10235
rect 13235 10199 13277 10523
rect 11983 10163 13277 10199
rect 11983 10129 11999 10163
rect 13075 10129 13091 10163
rect 11915 10101 11949 10117
rect 11915 9957 11949 9973
rect 13125 10101 13159 10117
rect 13125 9957 13159 9973
rect 10215 9914 11867 9931
rect 10537 9911 11867 9914
rect 11983 9911 11999 9945
rect 13075 9911 13091 9945
rect 10537 9899 13091 9911
rect 10537 9865 10553 9899
rect 11629 9897 13091 9899
rect 11629 9865 11645 9897
rect 11779 9875 13091 9897
rect 10469 9837 10503 9853
rect 10469 9653 10503 9669
rect 11679 9837 11713 9853
rect 11679 9653 11713 9669
rect 10537 9607 10553 9641
rect 11629 9607 11645 9641
rect 10365 9573 11645 9607
rect 10365 9307 10401 9573
rect 11779 9551 11839 9875
rect 13235 9839 13277 10163
rect 11983 9803 13277 9839
rect 11983 9769 11999 9803
rect 13075 9769 13091 9803
rect 11915 9741 11949 9757
rect 11915 9597 11949 9613
rect 13125 9741 13159 9757
rect 13125 9597 13159 9613
rect 11983 9551 11999 9585
rect 13075 9551 13091 9585
rect 11779 9515 13091 9551
rect 11779 9509 11839 9515
rect 10537 9475 11839 9509
rect 13235 9479 13277 9803
rect 10537 9441 10553 9475
rect 11629 9441 11645 9475
rect 10258 9291 10401 9307
rect 10376 9187 10401 9291
rect 10469 9413 10503 9429
rect 10469 9229 10503 9245
rect 11679 9413 11713 9429
rect 11679 9229 11713 9245
rect 10537 9187 10553 9217
rect 10376 9183 10553 9187
rect 11629 9183 11645 9217
rect 10376 9173 11645 9183
rect 10258 9158 11645 9173
rect 11797 9191 11839 9475
rect 11983 9443 13277 9479
rect 11983 9409 11999 9443
rect 13075 9409 13091 9443
rect 11915 9381 11949 9397
rect 11915 9237 11949 9253
rect 13125 9381 13159 9397
rect 13125 9237 13159 9253
rect 11983 9191 11999 9225
rect 13075 9191 13091 9225
rect 10258 9157 11575 9158
rect 10122 9128 10156 9154
rect 10365 9153 11575 9157
rect 11797 9155 13091 9191
rect 8861 9094 8921 9128
rect 9407 9094 9610 9128
rect 10096 9094 10156 9128
rect 7442 9056 8672 9061
rect 5718 8966 5734 9056
rect 8648 8966 8672 9056
rect 9467 9022 9550 9094
rect 10589 9061 11575 9153
rect 10345 9056 11575 9061
rect 8388 8961 8672 8966
rect 8861 8988 8921 9022
rect 9407 8988 9610 9022
rect 10096 8988 10156 9022
rect 8861 8962 8895 8988
rect 5740 8857 7034 8893
rect 5740 8533 5782 8857
rect 5926 8823 5942 8857
rect 7018 8823 7034 8857
rect 7400 8813 8861 8859
rect 5858 8795 5892 8811
rect 5858 8651 5892 8667
rect 7068 8795 7102 8811
rect 7402 8779 7418 8813
rect 8494 8779 8510 8813
rect 7334 8751 7368 8767
rect 7334 8687 7368 8703
rect 8544 8751 8578 8767
rect 8544 8687 8578 8703
rect 7068 8651 7102 8667
rect 7238 8645 7278 8673
rect 7402 8645 7418 8675
rect 7238 8641 7418 8645
rect 8494 8641 8510 8675
rect 5926 8605 5942 8639
rect 7018 8605 7034 8639
rect 7238 8605 7622 8641
rect 5926 8569 7186 8605
rect 5740 8497 7034 8533
rect 5740 8173 5782 8497
rect 5926 8463 5942 8497
rect 7018 8463 7034 8497
rect 5858 8435 5892 8451
rect 5858 8291 5892 8307
rect 7068 8435 7102 8451
rect 7068 8291 7102 8307
rect 5926 8245 5942 8279
rect 7018 8245 7034 8279
rect 7150 8265 7186 8569
rect 7238 8351 7278 8605
rect 8640 8555 8680 8813
rect 7400 8515 8680 8555
rect 7400 8509 7418 8515
rect 7402 8481 7418 8509
rect 8494 8509 8680 8515
rect 8494 8481 8510 8509
rect 8730 8498 8802 8522
rect 7334 8453 7368 8469
rect 7334 8389 7368 8405
rect 8544 8453 8578 8469
rect 8544 8389 8578 8405
rect 8730 8415 8748 8498
rect 8783 8415 8802 8498
rect 7402 8351 7418 8377
rect 7238 8343 7418 8351
rect 8494 8343 8510 8377
rect 7238 8309 7670 8343
rect 8730 8284 8802 8415
rect 8298 8265 8802 8284
rect 7150 8248 8802 8265
rect 7150 8245 8480 8248
rect 5926 8233 8480 8245
rect 5926 8231 7388 8233
rect 5926 8209 7238 8231
rect 5740 8137 7034 8173
rect 5740 7813 5782 8137
rect 5926 8103 5942 8137
rect 7018 8103 7034 8137
rect 5858 8075 5892 8091
rect 5858 7931 5892 7947
rect 7068 8075 7102 8091
rect 7068 7931 7102 7947
rect 5926 7885 5942 7919
rect 7018 7885 7034 7919
rect 7178 7885 7238 8209
rect 7372 8199 7388 8231
rect 8464 8199 8480 8233
rect 7304 8171 7338 8187
rect 7304 7987 7338 8003
rect 8514 8171 8548 8187
rect 8514 7987 8548 8003
rect 7372 7941 7388 7975
rect 8464 7941 8480 7975
rect 7372 7907 8652 7941
rect 5926 7849 7238 7885
rect 7178 7843 7238 7849
rect 5740 7777 7034 7813
rect 5926 7743 5942 7777
rect 7018 7743 7034 7777
rect 7178 7809 8480 7843
rect 5858 7715 5892 7731
rect 5858 7571 5892 7587
rect 7068 7715 7102 7731
rect 7068 7571 7102 7587
rect 5926 7525 5942 7559
rect 7018 7525 7034 7559
rect 7178 7525 7220 7809
rect 7372 7775 7388 7809
rect 8464 7775 8480 7809
rect 7304 7747 7338 7763
rect 7304 7563 7338 7579
rect 8514 7747 8548 7763
rect 8514 7563 8548 7579
rect 8616 7641 8652 7907
rect 8616 7625 8759 7641
rect 5926 7489 7220 7525
rect 7372 7517 7388 7551
rect 8464 7521 8480 7551
rect 8616 7521 8641 7625
rect 8464 7517 8641 7521
rect 7372 7507 8641 7517
rect 7372 7492 8759 7507
rect 7442 7491 8759 7492
rect 7442 7487 8652 7491
rect 9336 8962 9681 8988
rect 9336 8904 9433 8962
rect 9059 8854 9075 8888
rect 9251 8854 9267 8888
rect 8944 8826 9016 8842
rect 8944 8698 8982 8826
rect 8944 8682 9016 8698
rect 9310 8826 9381 8842
rect 9344 8698 9381 8826
rect 9310 8682 9381 8698
rect 8944 8556 8982 8682
rect 9059 8636 9075 8670
rect 9251 8636 9267 8670
rect 9344 8600 9381 8682
rect 9210 8578 9397 8600
rect 8944 8517 9115 8556
rect 9059 8480 9115 8517
rect 9210 8530 9274 8578
rect 9371 8530 9397 8578
rect 9210 8515 9397 8530
rect 9211 8480 9267 8515
rect 9059 8446 9075 8480
rect 9251 8446 9267 8480
rect 8982 8418 9016 8434
rect 8982 8164 9016 8290
rect 9310 8418 9344 8434
rect 9059 8228 9075 8262
rect 9251 8228 9267 8262
rect 9310 8187 9344 8290
rect 9271 8165 9376 8187
rect 9271 8164 9291 8165
rect 8982 8116 9291 8164
rect 8982 7972 9016 8116
rect 9271 8097 9291 8116
rect 9354 8097 9376 8165
rect 9271 8080 9376 8097
rect 9059 8000 9075 8034
rect 9251 8000 9267 8034
rect 8982 7588 9016 7604
rect 9310 7972 9344 8080
rect 9310 7588 9344 7604
rect 7442 7292 8428 7487
rect 8861 7462 8895 7488
rect 9058 7576 9268 7577
rect 9058 7542 9075 7576
rect 9251 7542 9268 7576
rect 9058 7462 9268 7542
rect 9467 7488 9550 8962
rect 9584 8904 9681 8962
rect 10122 8962 10156 8988
rect 9750 8854 9766 8888
rect 9942 8854 9958 8888
rect 9636 8826 9707 8842
rect 9636 8698 9673 8826
rect 9636 8682 9707 8698
rect 10001 8826 10073 8842
rect 10035 8698 10073 8826
rect 10001 8682 10073 8698
rect 9636 8600 9673 8682
rect 9750 8636 9766 8670
rect 9942 8636 9958 8670
rect 9620 8578 9807 8600
rect 9620 8530 9646 8578
rect 9743 8530 9807 8578
rect 10035 8556 10073 8682
rect 9620 8515 9807 8530
rect 9902 8517 10073 8556
rect 9750 8480 9806 8515
rect 9902 8480 9958 8517
rect 9750 8446 9766 8480
rect 9942 8446 9958 8480
rect 9673 8418 9707 8434
rect 9673 8187 9707 8290
rect 10001 8418 10035 8434
rect 9750 8228 9766 8262
rect 9942 8228 9958 8262
rect 9641 8165 9746 8187
rect 9641 8097 9663 8165
rect 9726 8164 9746 8165
rect 10001 8164 10035 8290
rect 9726 8116 10035 8164
rect 9726 8097 9746 8116
rect 9641 8080 9746 8097
rect 9673 7972 9707 8080
rect 9750 8000 9766 8034
rect 9942 8000 9958 8034
rect 9673 7588 9707 7604
rect 10001 7972 10035 8116
rect 10001 7588 10035 7604
rect 9433 7462 9584 7488
rect 9749 7576 9959 7577
rect 9749 7542 9766 7576
rect 9942 7542 9959 7576
rect 9749 7462 9959 7542
rect 10345 8966 10369 9056
rect 13283 8966 13299 9056
rect 10345 8961 10629 8966
rect 10156 8813 11617 8859
rect 11983 8857 13277 8893
rect 11983 8823 11999 8857
rect 13075 8823 13091 8857
rect 10337 8555 10377 8813
rect 10507 8779 10523 8813
rect 11599 8779 11615 8813
rect 11915 8795 11949 8811
rect 10439 8751 10473 8767
rect 10439 8687 10473 8703
rect 11649 8751 11683 8767
rect 11649 8687 11683 8703
rect 10507 8641 10523 8675
rect 11599 8645 11615 8675
rect 11739 8645 11779 8673
rect 11915 8651 11949 8667
rect 13125 8795 13159 8811
rect 13125 8651 13159 8667
rect 11599 8641 11779 8645
rect 11395 8605 11779 8641
rect 11983 8605 11999 8639
rect 13075 8605 13091 8639
rect 10215 8498 10287 8522
rect 10337 8515 11617 8555
rect 10337 8509 10523 8515
rect 10215 8415 10234 8498
rect 10269 8415 10287 8498
rect 10507 8481 10523 8509
rect 11599 8509 11617 8515
rect 11599 8481 11615 8509
rect 10215 8284 10287 8415
rect 10439 8453 10473 8469
rect 10439 8389 10473 8405
rect 11649 8453 11683 8469
rect 11649 8389 11683 8405
rect 10507 8343 10523 8377
rect 11599 8351 11615 8377
rect 11739 8351 11779 8605
rect 11599 8343 11779 8351
rect 11347 8309 11779 8343
rect 11831 8569 13091 8605
rect 10215 8265 10719 8284
rect 11831 8265 11867 8569
rect 13235 8533 13277 8857
rect 11983 8497 13277 8533
rect 11983 8463 11999 8497
rect 13075 8463 13091 8497
rect 11915 8435 11949 8451
rect 11915 8291 11949 8307
rect 13125 8435 13159 8451
rect 13125 8291 13159 8307
rect 10215 8248 11867 8265
rect 10537 8245 11867 8248
rect 11983 8245 11999 8279
rect 13075 8245 13091 8279
rect 10537 8233 13091 8245
rect 10537 8199 10553 8233
rect 11629 8231 13091 8233
rect 11629 8199 11645 8231
rect 11779 8209 13091 8231
rect 10469 8171 10503 8187
rect 10469 7987 10503 8003
rect 11679 8171 11713 8187
rect 11679 7987 11713 8003
rect 10537 7941 10553 7975
rect 11629 7941 11645 7975
rect 10365 7907 11645 7941
rect 10365 7641 10401 7907
rect 11779 7885 11839 8209
rect 13235 8173 13277 8497
rect 11983 8137 13277 8173
rect 11983 8103 11999 8137
rect 13075 8103 13091 8137
rect 11915 8075 11949 8091
rect 11915 7931 11949 7947
rect 13125 8075 13159 8091
rect 13125 7931 13159 7947
rect 11983 7885 11999 7919
rect 13075 7885 13091 7919
rect 11779 7849 13091 7885
rect 11779 7843 11839 7849
rect 10537 7809 11839 7843
rect 13235 7813 13277 8137
rect 10537 7775 10553 7809
rect 11629 7775 11645 7809
rect 10258 7625 10401 7641
rect 10376 7521 10401 7625
rect 10469 7747 10503 7763
rect 10469 7563 10503 7579
rect 11679 7747 11713 7763
rect 11679 7563 11713 7579
rect 10537 7521 10553 7551
rect 10376 7517 10553 7521
rect 11629 7517 11645 7551
rect 10376 7507 11645 7517
rect 10258 7492 11645 7507
rect 11797 7525 11839 7809
rect 11983 7777 13277 7813
rect 11983 7743 11999 7777
rect 13075 7743 13091 7777
rect 11915 7715 11949 7731
rect 11915 7571 11949 7587
rect 13125 7715 13159 7731
rect 13125 7571 13159 7587
rect 11983 7525 11999 7559
rect 13075 7525 13091 7559
rect 10258 7491 11575 7492
rect 10122 7462 10156 7488
rect 10365 7487 11575 7491
rect 11797 7489 13091 7525
rect 8861 7428 8921 7462
rect 9407 7428 9610 7462
rect 10096 7428 10156 7462
rect 10589 7292 11575 7487
rect 5606 7284 5735 7292
rect -1047 7076 2091 7226
rect 5452 7212 5735 7284
rect 13377 7284 13411 7292
rect 14530 18057 14644 18198
rect 18041 18198 18330 18214
rect 18041 18057 18152 18198
rect 14750 17836 14810 17870
rect 15463 17836 15523 17870
rect 14750 17810 14784 17836
rect 15489 17810 15523 17836
rect 15055 17732 15117 17766
rect 15155 17732 15217 17766
rect 15055 17673 15089 17732
rect 15055 15918 15089 15977
rect 15183 17673 15217 17732
rect 15183 15918 15217 15977
rect 15055 15884 15117 15918
rect 15155 15884 15217 15918
rect 14750 15823 14784 15849
rect 16247 17658 17282 18057
rect 15808 17618 15928 17658
rect 15523 17554 15664 17580
rect 15523 17386 15534 17554
rect 15635 17386 15664 17554
rect 15523 17362 15664 17386
rect 15882 17590 15928 17618
rect 17742 17618 17896 17658
rect 17742 17590 17822 17618
rect 16234 17462 16250 17496
rect 17426 17462 17442 17496
rect 16166 17434 16200 17450
rect 16166 17272 16200 17288
rect 17476 17434 17510 17450
rect 17476 17272 17510 17288
rect 16234 17226 16250 17260
rect 17426 17226 17442 17260
rect 16234 17092 16250 17126
rect 17426 17092 17442 17126
rect 16166 17064 16200 17080
rect 16166 16902 16200 16918
rect 17476 17064 17510 17080
rect 17476 16902 17510 16918
rect 16234 16856 16250 16890
rect 17426 16856 17442 16890
rect 16532 16694 16548 16728
rect 17136 16694 17152 16728
rect 16486 16644 16520 16660
rect 16486 16308 16520 16324
rect 17164 16644 17198 16660
rect 17420 16622 17436 16656
rect 17614 16622 17630 16656
rect 17374 16572 17408 16588
rect 17374 16416 17408 16432
rect 17642 16572 17822 16588
rect 17676 16432 17822 16572
rect 17642 16416 17822 16432
rect 17420 16348 17436 16382
rect 17614 16348 17630 16382
rect 17164 16308 17198 16324
rect 16532 16240 16548 16274
rect 17136 16240 17152 16274
rect 15882 16052 15954 16092
rect 15808 16024 15954 16052
rect 17648 16024 17724 16092
rect 17768 16052 17822 16092
rect 17768 16024 17896 16052
rect 15489 15823 15523 15849
rect 14750 15789 14810 15823
rect 15463 15789 15523 15823
rect 16361 15605 17268 16024
rect 14530 15597 18152 15605
rect 14530 15473 14634 15597
rect 14352 15440 14634 15473
rect 18031 15473 18152 15597
rect 18031 15440 18330 15473
rect 14387 13772 14444 13864
rect 18497 13772 18637 13864
rect 14387 13722 14466 13772
rect 18551 13756 18637 13772
rect 14764 13644 14824 13678
rect 17845 13660 17905 13678
rect 17845 13644 18317 13660
rect 14764 13618 18317 13644
rect 14798 13509 17871 13618
rect 14798 13456 14919 13509
rect 14978 13505 17871 13509
rect 14978 13502 17664 13505
rect 14978 13468 14994 13502
rect 15148 13468 15164 13502
rect 15478 13468 15494 13502
rect 15648 13468 15664 13502
rect 15978 13468 15994 13502
rect 16148 13468 16164 13502
rect 16478 13468 16494 13502
rect 16648 13468 16664 13502
rect 16978 13468 16994 13502
rect 17148 13468 17164 13502
rect 17478 13468 17494 13502
rect 17648 13468 17664 13502
rect 17720 13456 17871 13505
rect 14798 13440 14935 13456
rect 14798 12694 14901 13440
rect 14798 12678 14935 12694
rect 15207 13440 15241 13456
rect 15207 12678 15241 12694
rect 15401 13440 15435 13456
rect 15401 12678 15435 12694
rect 15707 13440 15741 13456
rect 15707 12678 15741 12694
rect 15901 13440 15935 13456
rect 15901 12678 15935 12694
rect 16207 13440 16241 13456
rect 16207 12678 16241 12694
rect 16401 13440 16435 13456
rect 16401 12678 16435 12694
rect 16707 13440 16741 13456
rect 16707 12678 16741 12694
rect 16901 13440 16935 13456
rect 16901 12678 16935 12694
rect 17207 13440 17241 13456
rect 17207 12678 17241 12694
rect 17401 13440 17435 13456
rect 17401 12678 17435 12694
rect 17707 13440 17871 13456
rect 17741 12694 17871 13440
rect 17707 12678 17871 12694
rect 14798 12517 14918 12678
rect 14978 12632 14994 12666
rect 15148 12632 15164 12666
rect 15478 12632 15494 12666
rect 15648 12632 15664 12666
rect 15978 12632 15994 12666
rect 16148 12632 16164 12666
rect 16478 12632 16494 12666
rect 16648 12632 16664 12666
rect 16978 12632 16994 12666
rect 17148 12632 17164 12666
rect 17478 12632 17494 12666
rect 17648 12632 17664 12666
rect 14764 12491 14918 12517
rect 15033 12491 15113 12632
rect 17536 12491 17616 12632
rect 17724 12517 17871 12678
rect 17905 13538 18317 13618
rect 17905 12517 18062 13538
rect 17724 12491 18062 12517
rect 14764 12457 14824 12491
rect 17845 12457 18062 12491
rect 14387 11848 14466 12335
rect 17626 12101 18062 12457
rect 18236 12101 18317 13538
rect 17626 11988 18317 12101
rect 14387 11838 14484 11848
rect 14299 11814 14484 11838
rect 14898 11814 14994 11848
rect 14299 11752 14422 11814
rect 14299 9302 14388 11752
rect 14960 11752 14994 11814
rect 14548 11712 14564 11746
rect 14818 11712 14834 11746
rect 14502 11662 14536 11678
rect 14502 10632 14536 10648
rect 14846 11662 14880 11678
rect 14846 10632 14880 10648
rect 14548 10564 14564 10598
rect 14818 10564 14834 10598
rect 14548 10456 14564 10490
rect 14818 10456 14834 10490
rect 14502 10406 14536 10422
rect 14502 9376 14536 9392
rect 14846 10406 14880 10422
rect 14846 9376 14880 9392
rect 14548 9308 14564 9342
rect 14818 9308 14834 9342
rect 14299 9240 14422 9302
rect 17626 11461 17892 11988
rect 16903 11427 16999 11461
rect 18207 11427 18303 11461
rect 16903 11365 16937 11427
rect 17478 11347 17762 11427
rect 18269 11365 18303 11427
rect 17082 11313 17098 11347
rect 18108 11313 18124 11347
rect 17005 11285 17039 11301
rect 17005 11227 17039 11243
rect 18167 11285 18201 11301
rect 18167 11227 18201 11243
rect 17082 11181 17098 11215
rect 18108 11181 18124 11215
rect 16903 11101 16937 11163
rect 18269 11101 18303 11163
rect 16903 11067 16999 11101
rect 18207 11067 18303 11101
rect 17481 10602 17709 10667
rect 17481 10441 17513 10602
rect 17670 10441 17709 10602
rect 14960 9240 14994 9302
rect 14299 9206 14484 9240
rect 14898 9206 14994 9240
rect 16843 10407 16903 10441
rect 18382 10407 18442 10441
rect 16843 10381 16877 10407
rect 17374 10323 17513 10407
rect 17670 10323 17849 10407
rect 17374 10280 17849 10323
rect 18408 10381 18442 10407
rect 17025 10246 17041 10280
rect 18231 10246 18247 10280
rect 16936 10218 16982 10234
rect 16936 9996 16948 10218
rect 16936 9618 16982 9996
rect 18290 10218 18336 10234
rect 18324 9996 18336 10218
rect 17025 9934 17041 9968
rect 18231 9934 18247 9968
rect 17025 9646 17041 9680
rect 18231 9646 18247 9680
rect 16936 9396 16948 9618
rect 16936 9380 16982 9396
rect 18290 9618 18336 9996
rect 18324 9396 18336 9618
rect 18290 9380 18336 9396
rect 17025 9334 17041 9368
rect 18231 9334 18247 9368
rect 14299 8850 14975 9206
rect 16843 9203 16877 9229
rect 18408 9203 18442 9229
rect 16843 9169 16903 9203
rect 18382 9169 18442 9203
rect 14298 8766 14383 8850
rect 18441 8842 18486 8850
rect 18441 8766 18551 8842
rect 14298 8693 14629 8766
rect 14380 8670 14629 8693
rect 14922 8670 17854 8704
rect 18148 8675 18551 8766
rect 18148 8670 18404 8675
rect 14380 8644 14538 8670
rect 14380 8602 14482 8644
rect 14522 8636 14538 8644
rect 14638 8636 14700 8670
rect 14922 8636 14938 8670
rect 15038 8636 15054 8670
rect 15322 8636 15338 8670
rect 15438 8636 15454 8670
rect 15722 8636 15738 8670
rect 15838 8636 15854 8670
rect 16122 8636 16138 8670
rect 16238 8636 16254 8670
rect 16522 8636 16538 8670
rect 16638 8636 16654 8670
rect 16922 8636 16938 8670
rect 17038 8636 17054 8670
rect 17322 8636 17338 8670
rect 17438 8636 17454 8670
rect 17722 8636 17738 8670
rect 17838 8636 17854 8670
rect 18076 8636 18138 8670
rect 18238 8636 18404 8670
rect 14654 8602 14700 8636
rect 18076 8602 18122 8636
rect 18285 8602 18404 8636
rect 14380 8586 14510 8602
rect 14380 7590 14476 8586
rect 14380 7574 14510 7590
rect 14666 8586 14700 8602
rect 14666 7574 14700 7590
rect 14831 8586 14910 8602
rect 14831 7590 14876 8586
rect 14831 7574 14910 7590
rect 15066 8586 15100 8602
rect 15066 7574 15100 7590
rect 15231 8586 15310 8602
rect 15231 7590 15276 8586
rect 15231 7574 15310 7590
rect 15466 8586 15500 8602
rect 15466 7574 15500 7590
rect 15631 8586 15710 8602
rect 15631 7590 15676 8586
rect 15631 7574 15710 7590
rect 15866 8586 15900 8602
rect 15866 7574 15900 7590
rect 16031 8586 16110 8602
rect 16031 7590 16076 8586
rect 16031 7574 16110 7590
rect 16266 8586 16300 8602
rect 16266 7574 16300 7590
rect 16476 8586 16510 8602
rect 16476 7574 16510 7590
rect 16666 8586 16745 8602
rect 16700 7590 16745 8586
rect 16666 7574 16745 7590
rect 16876 8586 16910 8602
rect 16876 7574 16910 7590
rect 17066 8586 17145 8602
rect 17100 7590 17145 8586
rect 17066 7574 17145 7590
rect 17276 8586 17310 8602
rect 17276 7574 17310 7590
rect 17466 8586 17545 8602
rect 17500 7590 17545 8586
rect 17466 7574 17545 7590
rect 17676 8586 17710 8602
rect 17676 7574 17710 7590
rect 17866 8586 17945 8602
rect 17900 7590 17945 8586
rect 17866 7574 17945 7590
rect 18076 8586 18110 8602
rect 18076 7574 18110 7590
rect 18266 8586 18404 8602
rect 18300 7590 18404 8586
rect 14380 7540 14482 7574
rect 14380 7529 14538 7540
rect 14298 7506 14538 7529
rect 14638 7506 14654 7540
rect 14298 7430 14631 7506
rect 14831 7430 14876 7574
rect 14922 7506 14938 7540
rect 15038 7506 15054 7540
rect 15231 7430 15276 7574
rect 15322 7506 15338 7540
rect 15438 7506 15454 7540
rect 15631 7430 15676 7574
rect 15722 7506 15738 7540
rect 15838 7506 15854 7540
rect 16031 7430 16076 7574
rect 16122 7506 16138 7540
rect 16238 7506 16254 7540
rect 16522 7506 16538 7540
rect 16638 7506 16654 7540
rect 16700 7430 16745 7574
rect 16922 7506 16938 7540
rect 17038 7506 17054 7540
rect 17100 7430 17145 7574
rect 17322 7506 17338 7540
rect 17438 7506 17454 7540
rect 17500 7430 17545 7574
rect 17722 7506 17738 7540
rect 17838 7506 17854 7540
rect 17900 7430 17945 7574
rect 18266 7540 18404 7590
rect 18122 7506 18138 7540
rect 18238 7511 18404 7540
rect 18486 7511 18551 8675
rect 18238 7506 18551 7511
rect 18146 7430 18551 7506
rect 14298 7386 14383 7430
rect 13377 7212 13565 7284
rect 14296 7346 14383 7386
rect 18441 7350 18551 7430
rect 18441 7346 18637 7350
rect 5959 7076 12804 7212
rect 14296 7076 15868 7346
rect 18155 7327 18637 7346
rect 18155 7076 18635 7327
rect -1047 6476 18788 7076
rect -1047 6466 -494 6476
<< viali >>
rect -69 18995 407 19029
rect -153 18799 -119 18967
rect 457 18799 491 18967
rect -69 18737 407 18771
rect -69 18579 407 18613
rect -153 18383 -119 18551
rect 457 18383 491 18551
rect -69 18321 407 18355
rect -69 18163 407 18197
rect -153 17967 -119 18135
rect 457 17967 491 18135
rect -69 17905 407 17939
rect -69 17747 407 17781
rect -153 17551 -119 17719
rect 457 17551 491 17719
rect -69 17489 407 17523
rect -69 17331 407 17365
rect -153 17135 -119 17303
rect 457 17135 491 17303
rect -69 17073 407 17107
rect -69 16915 407 16949
rect -153 16719 -119 16887
rect 457 16719 491 16887
rect -69 16657 407 16691
rect -69 16499 407 16533
rect -153 16303 -119 16471
rect 457 16303 491 16471
rect -69 16241 407 16275
rect -69 16083 407 16117
rect -153 15887 -119 16055
rect 457 15887 491 16055
rect -69 15825 407 15859
rect 1402 19245 1770 19279
rect 1340 19110 1374 19186
rect 1798 19110 1832 19186
rect 1402 19017 1770 19051
rect 2102 19245 2470 19279
rect 2040 19110 2074 19186
rect 2498 19110 2532 19186
rect 2102 19017 2470 19051
rect 1402 18861 1770 18895
rect 2102 18861 2470 18895
rect 1340 18326 1374 18802
rect 1798 18326 1832 18802
rect 1898 18539 1954 18603
rect 2040 18326 2074 18802
rect 2498 18326 2532 18802
rect 1402 18233 1770 18267
rect 2102 18233 2470 18267
rect 1402 18077 1770 18111
rect 2102 18077 2470 18111
rect 1340 17542 1374 18018
rect 1798 17542 1832 18018
rect 1402 17449 1770 17483
rect 1402 17293 1770 17327
rect 1340 16758 1374 17234
rect 1798 16758 1832 17234
rect 2040 17542 2074 18018
rect 2498 17542 2532 18018
rect 2102 17449 2470 17483
rect 2102 17293 2470 17327
rect 2040 16758 2074 17234
rect 2498 16758 2532 17234
rect 1402 16665 1770 16699
rect 2102 16665 2470 16699
rect 1402 16509 1770 16543
rect 2102 16509 2470 16543
rect 1340 15974 1374 16450
rect 1798 15974 1832 16450
rect 1901 16177 1957 16241
rect 2040 15974 2074 16450
rect 2498 15974 2532 16450
rect 1167 15765 1256 15945
rect 1402 15881 1770 15915
rect 2102 15881 2470 15915
rect 1402 15725 1770 15759
rect 1340 15590 1374 15666
rect 1798 15590 1832 15666
rect 1402 15497 1770 15531
rect 2102 15725 2470 15759
rect 2040 15590 2074 15666
rect 2498 15590 2532 15666
rect 2102 15497 2470 15531
rect 70 14651 238 14685
rect 486 14651 654 14685
rect 902 14651 1070 14685
rect 1318 14651 1486 14685
rect 1734 14651 1902 14685
rect 2150 14651 2318 14685
rect 8 14125 42 14601
rect 266 14125 300 14601
rect 70 14041 238 14075
rect 424 14125 458 14601
rect 682 14125 716 14601
rect 840 14125 874 14601
rect 1098 14125 1132 14601
rect 1256 14125 1290 14601
rect 1514 14125 1548 14601
rect 1672 14125 1706 14601
rect 1930 14125 1964 14601
rect 2088 14125 2122 14601
rect 2346 14125 2380 14601
rect 486 14041 654 14075
rect 902 14041 1070 14075
rect 1318 14041 1486 14075
rect 964 13946 1084 13983
rect 1734 14041 1902 14075
rect 2150 14041 2318 14075
rect 675 13767 1643 13801
rect 613 13541 647 13717
rect 1671 13541 1705 13717
rect 675 13457 1643 13491
rect 1185 13005 1366 13218
rect -151 12692 225 12726
rect 485 12692 861 12726
rect 1121 12692 1497 12726
rect 1757 12692 2133 12726
rect -244 12596 -210 12664
rect 284 12596 318 12664
rect 392 12596 426 12664
rect 920 12596 954 12664
rect 1028 12596 1062 12664
rect 1556 12596 1590 12664
rect 1664 12596 1698 12664
rect 2192 12596 2226 12664
rect -151 12534 225 12568
rect 485 12534 861 12568
rect 1121 12534 1497 12568
rect 1757 12534 2133 12568
rect 62 12308 146 12409
rect 2207 12260 2467 12331
rect 2467 12260 2491 12331
rect 795 11946 2157 11980
rect 733 11735 767 11887
rect 2185 11735 2219 11887
rect 795 11642 2157 11676
rect 698 11357 875 11510
rect 417 11044 939 11078
rect 355 10323 389 10985
rect 967 10323 1001 10985
rect 417 10230 939 10264
rect 1411 11038 2179 11072
rect 1349 10903 1383 10979
rect 2207 10903 2241 10979
rect 1411 10810 2179 10844
rect 1337 10646 2181 10680
rect 1275 10137 1309 10587
rect 2209 10137 2243 10587
rect 1337 10044 2181 10078
rect 1171 9299 1539 9333
rect 1871 9299 2239 9333
rect 1109 8764 1143 9240
rect 1567 8764 1601 9240
rect 1809 8764 1843 9240
rect 2267 8764 2301 9240
rect 1171 8671 1539 8705
rect 1871 8671 2239 8705
rect 1171 8515 1539 8549
rect 1871 8515 2239 8549
rect 2420 8504 2433 9116
rect 2433 8504 2762 9116
rect 1109 7980 1143 8456
rect 1567 7980 1601 8456
rect 1809 7980 1843 8456
rect 2267 7980 2301 8456
rect 1171 7887 1539 7921
rect 1871 7887 2239 7921
rect 3098 19261 3466 19295
rect 3036 19126 3070 19202
rect 3494 19126 3528 19202
rect 3798 19261 4166 19295
rect 3736 19126 3770 19202
rect 4194 19126 4228 19202
rect 3098 19033 3466 19067
rect 3798 19033 4166 19067
rect 3098 18877 3466 18911
rect 3798 18877 4166 18911
rect 3036 18342 3070 18818
rect 3494 18342 3528 18818
rect 3736 18342 3770 18818
rect 4194 18342 4228 18818
rect 3098 18249 3466 18283
rect 3798 18249 4166 18283
rect 3098 18093 3466 18127
rect 3798 18093 4166 18127
rect 3036 17558 3070 18034
rect 3494 17558 3528 18034
rect 3736 17558 3770 18034
rect 4194 17558 4228 18034
rect 3098 17465 3466 17499
rect 3798 17465 4166 17499
rect 3098 17309 3466 17343
rect 3798 17309 4166 17343
rect 3036 16774 3070 17250
rect 3494 16774 3528 17250
rect 3736 16774 3770 17250
rect 4194 16774 4228 17250
rect 3098 16681 3466 16715
rect 3798 16681 4166 16715
rect 3098 16525 3466 16559
rect 3798 16525 4166 16559
rect 3036 15990 3070 16466
rect 3494 15990 3528 16466
rect 3736 15990 3770 16466
rect 4194 15990 4228 16466
rect 3098 15897 3466 15931
rect 3798 15897 4166 15931
rect 3098 15741 3466 15775
rect 3798 15741 4166 15775
rect 3036 15206 3070 15682
rect 3494 15206 3528 15682
rect 3736 15206 3770 15682
rect 4194 15206 4228 15682
rect 3098 15113 3466 15147
rect 3798 15113 4166 15147
rect 3098 14957 3466 14991
rect 3798 14957 4166 14991
rect 3036 14422 3070 14898
rect 3494 14422 3528 14898
rect 3594 14635 3650 14699
rect 3736 14422 3770 14898
rect 4194 14422 4228 14898
rect 3098 14329 3466 14363
rect 3798 14329 4166 14363
rect 3098 14173 3466 14207
rect 3798 14173 4166 14207
rect 3036 13638 3070 14114
rect 3494 13638 3528 14114
rect 3098 13545 3466 13579
rect 3098 13389 3466 13423
rect 3036 12854 3070 13330
rect 3494 12854 3528 13330
rect 3736 13638 3770 14114
rect 4194 13638 4228 14114
rect 3798 13545 4166 13579
rect 3798 13389 4166 13423
rect 3736 12854 3770 13330
rect 4194 12854 4228 13330
rect 3098 12761 3466 12795
rect 3798 12761 4166 12795
rect 3098 12605 3466 12639
rect 3798 12605 4166 12639
rect 3036 12070 3070 12546
rect 3494 12070 3528 12546
rect 3597 12273 3653 12337
rect 3736 12070 3770 12546
rect 4194 12070 4228 12546
rect 3098 11977 3466 12011
rect 3798 11977 4166 12011
rect 3098 11821 3466 11855
rect 3798 11821 4166 11855
rect 3036 11286 3070 11762
rect 3494 11286 3528 11762
rect 3736 11286 3770 11762
rect 4194 11286 4228 11762
rect 3098 11193 3466 11227
rect 3798 11193 4166 11227
rect 3098 11037 3466 11071
rect 3798 11037 4166 11071
rect 3036 10502 3070 10978
rect 3494 10502 3528 10978
rect 3736 10502 3770 10978
rect 4194 10502 4228 10978
rect 3098 10409 3466 10443
rect 3798 10409 4166 10443
rect 3098 10253 3466 10287
rect 3798 10253 4166 10287
rect 3036 9718 3070 10194
rect 3494 9718 3528 10194
rect 3736 9718 3770 10194
rect 4194 9718 4228 10194
rect 3098 9625 3466 9659
rect 3798 9625 4166 9659
rect 3098 9469 3466 9503
rect 3798 9469 4166 9503
rect 3036 8934 3070 9410
rect 3494 8934 3528 9410
rect 3736 8934 3770 9410
rect 4194 8934 4228 9410
rect 3098 8841 3466 8875
rect 3798 8841 4166 8875
rect 3098 8685 3466 8719
rect 3798 8685 4166 8719
rect 3036 8150 3070 8626
rect 3494 8150 3528 8626
rect 3736 8150 3770 8626
rect 4194 8150 4228 8626
rect 3098 8057 3466 8091
rect 3798 8057 4166 8091
rect 3098 7901 3466 7935
rect 3798 7901 4166 7935
rect 3036 7766 3070 7842
rect 3494 7766 3528 7842
rect 3098 7673 3466 7707
rect 3736 7766 3770 7842
rect 4194 7766 4228 7842
rect 3798 7673 4166 7707
rect 7113 19565 10289 19644
rect 7113 19508 10289 19565
rect 5907 19305 6035 19339
rect 6307 19305 6435 19339
rect 6707 19305 6835 19339
rect 7107 19305 7235 19339
rect 7507 19305 7635 19339
rect 7907 19305 8035 19339
rect 8307 19305 8435 19339
rect 8707 19305 8835 19339
rect 9107 19305 9235 19339
rect 9507 19305 9635 19339
rect 9907 19305 10035 19339
rect 10307 19305 10435 19339
rect 10707 19305 10835 19339
rect 11107 19305 11235 19339
rect 11507 19305 11635 19339
rect 11907 19305 12035 19339
rect 5845 18179 5879 19255
rect 6063 18179 6097 19255
rect 6245 18179 6279 19255
rect 6463 18179 6497 19255
rect 6645 18179 6679 19255
rect 6863 18179 6897 19255
rect 7045 18179 7079 19255
rect 7263 18179 7297 19255
rect 7445 18179 7479 19255
rect 7663 18179 7697 19255
rect 7845 18179 7879 19255
rect 8063 18179 8097 19255
rect 8245 18179 8279 19255
rect 8463 18179 8497 19255
rect 8645 18179 8679 19255
rect 8863 18179 8897 19255
rect 9045 18179 9079 19255
rect 9263 18179 9297 19255
rect 9445 18179 9479 19255
rect 9663 18179 9697 19255
rect 9845 18179 9879 19255
rect 10063 18179 10097 19255
rect 10245 18179 10279 19255
rect 10463 18179 10497 19255
rect 10645 18179 10679 19255
rect 10863 18179 10897 19255
rect 11045 18179 11079 19255
rect 11263 18179 11297 19255
rect 11445 18179 11479 19255
rect 11663 18179 11697 19255
rect 11845 18179 11879 19255
rect 12063 18179 12097 19255
rect 5907 18095 6035 18129
rect 6307 18095 6435 18129
rect 6707 18095 6835 18129
rect 7107 18095 7235 18129
rect 7507 18095 7635 18129
rect 7907 18095 8035 18129
rect 8307 18095 8435 18129
rect 8707 18095 8835 18129
rect 9107 18095 9235 18129
rect 9507 18095 9635 18129
rect 9907 18095 10035 18129
rect 10307 18095 10435 18129
rect 10707 18095 10835 18129
rect 11107 18095 11235 18129
rect 11507 18095 11635 18129
rect 11907 18095 12035 18129
rect 10110 17718 10525 17815
rect 5786 17605 5914 17639
rect 6186 17605 6314 17639
rect 6586 17605 6714 17639
rect 6986 17605 7114 17639
rect 7386 17605 7514 17639
rect 7786 17605 7914 17639
rect 8186 17605 8314 17639
rect 8586 17605 8714 17639
rect 5724 16479 5758 17555
rect 5942 16479 5976 17555
rect 6124 16479 6158 17555
rect 6342 16479 6376 17555
rect 6524 16479 6558 17555
rect 6742 16479 6776 17555
rect 6924 16479 6958 17555
rect 7142 16479 7176 17555
rect 7324 16479 7358 17555
rect 7542 16479 7576 17555
rect 7724 16479 7758 17555
rect 7942 16479 7976 17555
rect 8124 16479 8158 17555
rect 8342 16479 8376 17555
rect 8524 16479 8558 17555
rect 8742 16479 8776 17555
rect 5786 16395 5914 16429
rect 6186 16395 6314 16429
rect 6586 16395 6714 16429
rect 6986 16395 7114 16429
rect 7386 16395 7514 16429
rect 7786 16395 7914 16429
rect 8186 16395 8314 16429
rect 8586 16395 8714 16429
rect 9430 17361 9558 17395
rect 9830 17361 9958 17395
rect 9368 17126 9402 17302
rect 9586 17126 9620 17302
rect 9768 17126 9802 17302
rect 9430 17033 9558 17067
rect 9986 17126 10020 17302
rect 9830 17033 9958 17067
rect 10689 17332 10817 17366
rect 11089 17332 11217 17366
rect 11489 17332 11617 17366
rect 11889 17332 12017 17366
rect 10627 17097 10661 17273
rect 10845 17097 10879 17273
rect 11027 17097 11061 17273
rect 11245 17097 11279 17273
rect 11427 17097 11461 17273
rect 11645 17097 11679 17273
rect 11827 17097 11861 17273
rect 12045 17097 12079 17273
rect 10689 17004 10817 17038
rect 11089 17004 11217 17038
rect 11489 17004 11617 17038
rect 11889 17004 12017 17038
rect 11180 16762 11520 16851
rect 9052 16375 9594 16473
rect 10546 16377 10771 16692
rect 6477 16165 7983 16264
rect 8416 15638 8643 15707
rect 9383 15686 9629 15974
rect 9383 15652 9407 15686
rect 9407 15652 9610 15686
rect 9610 15652 9629 15686
rect 5942 15487 7018 15521
rect 5858 15331 5892 15459
rect 7068 15331 7102 15459
rect 7418 15443 8494 15477
rect 7334 15367 7368 15415
rect 8544 15367 8578 15415
rect 7418 15305 8494 15339
rect 5942 15269 7018 15303
rect 5942 15127 7018 15161
rect 5858 14971 5892 15099
rect 7068 14971 7102 15099
rect 5942 14909 7018 14943
rect 7418 15145 8494 15179
rect 7334 15069 7368 15117
rect 8544 15069 8578 15117
rect 8748 15079 8783 15162
rect 7418 15007 8494 15041
rect 5942 14767 7018 14801
rect 5858 14611 5892 14739
rect 7068 14611 7102 14739
rect 5942 14549 7018 14583
rect 7388 14863 8464 14897
rect 7304 14667 7338 14835
rect 8514 14667 8548 14835
rect 7388 14605 8464 14639
rect 5942 14407 7018 14441
rect 5858 14251 5892 14379
rect 7068 14251 7102 14379
rect 5942 14189 7018 14223
rect 7388 14439 8464 14473
rect 7304 14243 7338 14411
rect 8514 14243 8548 14411
rect 7388 14181 8464 14215
rect 9383 15626 9629 15652
rect 9383 15598 9433 15626
rect 9433 15598 9467 15626
rect 9467 15598 9550 15626
rect 9550 15598 9584 15626
rect 9584 15598 9629 15626
rect 9075 15518 9251 15552
rect 8982 15362 9016 15490
rect 9310 15362 9344 15490
rect 9075 15300 9251 15334
rect 9274 15194 9371 15242
rect 9075 15110 9251 15144
rect 8982 14954 9016 15082
rect 9310 14954 9344 15082
rect 9075 14892 9251 14926
rect 9291 14761 9354 14829
rect 9075 14664 9251 14698
rect 8982 14268 9016 14636
rect 9310 14268 9344 14636
rect 9075 14206 9251 14240
rect 9766 15518 9942 15552
rect 9673 15362 9707 15490
rect 10001 15362 10035 15490
rect 9766 15300 9942 15334
rect 9646 15194 9743 15242
rect 9766 15110 9942 15144
rect 9673 14954 9707 15082
rect 10001 14954 10035 15082
rect 9766 14892 9942 14926
rect 9663 14761 9726 14829
rect 9766 14664 9942 14698
rect 9673 14268 9707 14636
rect 10001 14268 10035 14636
rect 9766 14206 9942 14240
rect 10374 15638 10601 15707
rect 11999 15487 13075 15521
rect 10523 15443 11599 15477
rect 10439 15367 10473 15415
rect 11649 15367 11683 15415
rect 10523 15305 11599 15339
rect 11915 15331 11949 15459
rect 13125 15331 13159 15459
rect 11999 15269 13075 15303
rect 10234 15079 10269 15162
rect 10523 15145 11599 15179
rect 10439 15069 10473 15117
rect 11649 15069 11683 15117
rect 10523 15007 11599 15041
rect 11999 15127 13075 15161
rect 11915 14971 11949 15099
rect 13125 14971 13159 15099
rect 11999 14909 13075 14943
rect 10553 14863 11629 14897
rect 10469 14667 10503 14835
rect 11679 14667 11713 14835
rect 10553 14605 11629 14639
rect 11999 14767 13075 14801
rect 11915 14611 11949 14739
rect 13125 14611 13159 14739
rect 11999 14549 13075 14583
rect 10553 14439 11629 14473
rect 10469 14243 10503 14411
rect 11679 14243 11713 14411
rect 10553 14181 11629 14215
rect 11999 14407 13075 14441
rect 11915 14251 11949 14379
rect 13125 14251 13159 14379
rect 11999 14189 13075 14223
rect 8416 13972 8643 14041
rect 5942 13821 7018 13855
rect 5858 13665 5892 13793
rect 7068 13665 7102 13793
rect 7418 13777 8494 13811
rect 7334 13701 7368 13749
rect 8544 13701 8578 13749
rect 7418 13639 8494 13673
rect 5942 13603 7018 13637
rect 5942 13461 7018 13495
rect 5858 13305 5892 13433
rect 7068 13305 7102 13433
rect 5942 13243 7018 13277
rect 7418 13479 8494 13513
rect 7334 13403 7368 13451
rect 8544 13403 8578 13451
rect 8748 13413 8783 13496
rect 7418 13341 8494 13375
rect 5942 13101 7018 13135
rect 5858 12945 5892 13073
rect 7068 12945 7102 13073
rect 5942 12883 7018 12917
rect 7388 13197 8464 13231
rect 7304 13001 7338 13169
rect 8514 13001 8548 13169
rect 7388 12939 8464 12973
rect 5942 12741 7018 12775
rect 5858 12585 5892 12713
rect 7068 12585 7102 12713
rect 5942 12523 7018 12557
rect 7388 12773 8464 12807
rect 7304 12577 7338 12745
rect 8514 12577 8548 12745
rect 7388 12515 8464 12549
rect 9075 13852 9251 13886
rect 8982 13696 9016 13824
rect 9310 13696 9344 13824
rect 9075 13634 9251 13668
rect 9274 13528 9371 13576
rect 9075 13444 9251 13478
rect 8982 13288 9016 13416
rect 9310 13288 9344 13416
rect 9075 13226 9251 13260
rect 9291 13095 9354 13163
rect 9075 12998 9251 13032
rect 8982 12602 9016 12970
rect 9310 12602 9344 12970
rect 9075 12540 9251 12574
rect 9766 13852 9942 13886
rect 9673 13696 9707 13824
rect 10001 13696 10035 13824
rect 9766 13634 9942 13668
rect 9646 13528 9743 13576
rect 9766 13444 9942 13478
rect 9673 13288 9707 13416
rect 10001 13288 10035 13416
rect 9766 13226 9942 13260
rect 9663 13095 9726 13163
rect 9766 12998 9942 13032
rect 9673 12602 9707 12970
rect 10001 12602 10035 12970
rect 9766 12540 9942 12574
rect 10374 13972 10601 14041
rect 11999 13821 13075 13855
rect 10523 13777 11599 13811
rect 10439 13701 10473 13749
rect 11649 13701 11683 13749
rect 10523 13639 11599 13673
rect 11915 13665 11949 13793
rect 13125 13665 13159 13793
rect 11999 13603 13075 13637
rect 10234 13413 10269 13496
rect 10523 13479 11599 13513
rect 10439 13403 10473 13451
rect 11649 13403 11683 13451
rect 10523 13341 11599 13375
rect 11999 13461 13075 13495
rect 11915 13305 11949 13433
rect 13125 13305 13159 13433
rect 11999 13243 13075 13277
rect 10553 13197 11629 13231
rect 10469 13001 10503 13169
rect 11679 13001 11713 13169
rect 10553 12939 11629 12973
rect 11999 13101 13075 13135
rect 11915 12945 11949 13073
rect 13125 12945 13159 13073
rect 11999 12883 13075 12917
rect 10553 12773 11629 12807
rect 10469 12577 10503 12745
rect 11679 12577 11713 12745
rect 10553 12515 11629 12549
rect 11999 12741 13075 12775
rect 11915 12585 11949 12713
rect 13125 12585 13159 12713
rect 11999 12523 13075 12557
rect 8416 12306 8643 12375
rect 5942 12155 7018 12189
rect 5858 11999 5892 12127
rect 7068 11999 7102 12127
rect 7418 12111 8494 12145
rect 7334 12035 7368 12083
rect 8544 12035 8578 12083
rect 7418 11973 8494 12007
rect 5942 11937 7018 11971
rect 5942 11795 7018 11829
rect 5858 11639 5892 11767
rect 7068 11639 7102 11767
rect 5942 11577 7018 11611
rect 7418 11813 8494 11847
rect 7334 11737 7368 11785
rect 8544 11737 8578 11785
rect 8748 11747 8783 11830
rect 7418 11675 8494 11709
rect 5942 11435 7018 11469
rect 5858 11279 5892 11407
rect 7068 11279 7102 11407
rect 5942 11217 7018 11251
rect 7388 11531 8464 11565
rect 7304 11335 7338 11503
rect 8514 11335 8548 11503
rect 7388 11273 8464 11307
rect 5942 11075 7018 11109
rect 5858 10919 5892 11047
rect 7068 10919 7102 11047
rect 5942 10857 7018 10891
rect 7388 11107 8464 11141
rect 7304 10911 7338 11079
rect 8514 10911 8548 11079
rect 7388 10849 8464 10883
rect 9075 12186 9251 12220
rect 8982 12030 9016 12158
rect 9310 12030 9344 12158
rect 9075 11968 9251 12002
rect 9274 11862 9371 11910
rect 9075 11778 9251 11812
rect 8982 11622 9016 11750
rect 9310 11622 9344 11750
rect 9075 11560 9251 11594
rect 9291 11429 9354 11497
rect 9075 11332 9251 11366
rect 8982 10936 9016 11304
rect 9310 10936 9344 11304
rect 9075 10874 9251 10908
rect 9766 12186 9942 12220
rect 9673 12030 9707 12158
rect 10001 12030 10035 12158
rect 9766 11968 9942 12002
rect 9646 11862 9743 11910
rect 9766 11778 9942 11812
rect 9673 11622 9707 11750
rect 10001 11622 10035 11750
rect 9766 11560 9942 11594
rect 9663 11429 9726 11497
rect 9766 11332 9942 11366
rect 9673 10936 9707 11304
rect 10001 10936 10035 11304
rect 9766 10874 9942 10908
rect 10374 12306 10601 12375
rect 11999 12155 13075 12189
rect 10523 12111 11599 12145
rect 10439 12035 10473 12083
rect 11649 12035 11683 12083
rect 10523 11973 11599 12007
rect 11915 11999 11949 12127
rect 13125 11999 13159 12127
rect 11999 11937 13075 11971
rect 10234 11747 10269 11830
rect 10523 11813 11599 11847
rect 10439 11737 10473 11785
rect 11649 11737 11683 11785
rect 10523 11675 11599 11709
rect 11999 11795 13075 11829
rect 11915 11639 11949 11767
rect 13125 11639 13159 11767
rect 11999 11577 13075 11611
rect 10553 11531 11629 11565
rect 10469 11335 10503 11503
rect 11679 11335 11713 11503
rect 10553 11273 11629 11307
rect 11999 11435 13075 11469
rect 11915 11279 11949 11407
rect 13125 11279 13159 11407
rect 11999 11217 13075 11251
rect 10553 11107 11629 11141
rect 10469 10911 10503 11079
rect 11679 10911 11713 11079
rect 10553 10849 11629 10883
rect 11999 11075 13075 11109
rect 11915 10919 11949 11047
rect 13125 10919 13159 11047
rect 11999 10857 13075 10891
rect 8416 10640 8643 10709
rect 5942 10489 7018 10523
rect 5858 10333 5892 10461
rect 7068 10333 7102 10461
rect 7418 10445 8494 10479
rect 7334 10369 7368 10417
rect 8544 10369 8578 10417
rect 7418 10307 8494 10341
rect 5942 10271 7018 10305
rect 5942 10129 7018 10163
rect 5858 9973 5892 10101
rect 7068 9973 7102 10101
rect 5942 9911 7018 9945
rect 7418 10147 8494 10181
rect 7334 10071 7368 10119
rect 8544 10071 8578 10119
rect 8748 10081 8783 10164
rect 7418 10009 8494 10043
rect 5942 9769 7018 9803
rect 5858 9613 5892 9741
rect 7068 9613 7102 9741
rect 5942 9551 7018 9585
rect 7388 9865 8464 9899
rect 7304 9669 7338 9837
rect 8514 9669 8548 9837
rect 7388 9607 8464 9641
rect 5942 9409 7018 9443
rect 5858 9253 5892 9381
rect 7068 9253 7102 9381
rect 5942 9191 7018 9225
rect 7388 9441 8464 9475
rect 7304 9245 7338 9413
rect 8514 9245 8548 9413
rect 7388 9183 8464 9217
rect 9075 10520 9251 10554
rect 8982 10364 9016 10492
rect 9310 10364 9344 10492
rect 9075 10302 9251 10336
rect 9274 10196 9371 10244
rect 9075 10112 9251 10146
rect 8982 9956 9016 10084
rect 9310 9956 9344 10084
rect 9075 9894 9251 9928
rect 9291 9763 9354 9831
rect 9075 9666 9251 9700
rect 8982 9270 9016 9638
rect 9310 9270 9344 9638
rect 9075 9208 9251 9242
rect 9766 10520 9942 10554
rect 9673 10364 9707 10492
rect 10001 10364 10035 10492
rect 9766 10302 9942 10336
rect 9646 10196 9743 10244
rect 9766 10112 9942 10146
rect 9673 9956 9707 10084
rect 10001 9956 10035 10084
rect 9766 9894 9942 9928
rect 9663 9763 9726 9831
rect 9766 9666 9942 9700
rect 9673 9270 9707 9638
rect 10001 9270 10035 9638
rect 9766 9208 9942 9242
rect 10374 10640 10601 10709
rect 11999 10489 13075 10523
rect 10523 10445 11599 10479
rect 10439 10369 10473 10417
rect 11649 10369 11683 10417
rect 10523 10307 11599 10341
rect 11915 10333 11949 10461
rect 13125 10333 13159 10461
rect 11999 10271 13075 10305
rect 10234 10081 10269 10164
rect 10523 10147 11599 10181
rect 10439 10071 10473 10119
rect 11649 10071 11683 10119
rect 10523 10009 11599 10043
rect 11999 10129 13075 10163
rect 11915 9973 11949 10101
rect 13125 9973 13159 10101
rect 11999 9911 13075 9945
rect 10553 9865 11629 9899
rect 10469 9669 10503 9837
rect 11679 9669 11713 9837
rect 10553 9607 11629 9641
rect 11999 9769 13075 9803
rect 11915 9613 11949 9741
rect 13125 9613 13159 9741
rect 11999 9551 13075 9585
rect 10553 9441 11629 9475
rect 10469 9245 10503 9413
rect 11679 9245 11713 9413
rect 10553 9183 11629 9217
rect 11999 9409 13075 9443
rect 11915 9253 11949 9381
rect 13125 9253 13159 9381
rect 11999 9191 13075 9225
rect 8416 8974 8643 9043
rect 5942 8823 7018 8857
rect 5858 8667 5892 8795
rect 7068 8667 7102 8795
rect 7418 8779 8494 8813
rect 7334 8703 7368 8751
rect 8544 8703 8578 8751
rect 7418 8641 8494 8675
rect 5942 8605 7018 8639
rect 5942 8463 7018 8497
rect 5858 8307 5892 8435
rect 7068 8307 7102 8435
rect 5942 8245 7018 8279
rect 7418 8481 8494 8515
rect 7334 8405 7368 8453
rect 8544 8405 8578 8453
rect 8748 8415 8783 8498
rect 7418 8343 8494 8377
rect 5942 8103 7018 8137
rect 5858 7947 5892 8075
rect 7068 7947 7102 8075
rect 5942 7885 7018 7919
rect 7388 8199 8464 8233
rect 7304 8003 7338 8171
rect 8514 8003 8548 8171
rect 7388 7941 8464 7975
rect 5942 7743 7018 7777
rect 5858 7587 5892 7715
rect 7068 7587 7102 7715
rect 5942 7525 7018 7559
rect 7388 7775 8464 7809
rect 7304 7579 7338 7747
rect 8514 7579 8548 7747
rect 7388 7517 8464 7551
rect 9075 8854 9251 8888
rect 8982 8698 9016 8826
rect 9310 8698 9344 8826
rect 9075 8636 9251 8670
rect 9274 8530 9371 8578
rect 9075 8446 9251 8480
rect 8982 8290 9016 8418
rect 9310 8290 9344 8418
rect 9075 8228 9251 8262
rect 9291 8097 9354 8165
rect 9075 8000 9251 8034
rect 8982 7604 9016 7972
rect 9310 7604 9344 7972
rect 9075 7542 9251 7576
rect 9766 8854 9942 8888
rect 9673 8698 9707 8826
rect 10001 8698 10035 8826
rect 9766 8636 9942 8670
rect 9646 8530 9743 8578
rect 9766 8446 9942 8480
rect 9673 8290 9707 8418
rect 10001 8290 10035 8418
rect 9766 8228 9942 8262
rect 9663 8097 9726 8165
rect 9766 8000 9942 8034
rect 9673 7604 9707 7972
rect 10001 7604 10035 7972
rect 9766 7542 9942 7576
rect 10374 8974 10601 9043
rect 11999 8823 13075 8857
rect 10523 8779 11599 8813
rect 10439 8703 10473 8751
rect 11649 8703 11683 8751
rect 10523 8641 11599 8675
rect 11915 8667 11949 8795
rect 13125 8667 13159 8795
rect 11999 8605 13075 8639
rect 10234 8415 10269 8498
rect 10523 8481 11599 8515
rect 10439 8405 10473 8453
rect 11649 8405 11683 8453
rect 10523 8343 11599 8377
rect 11999 8463 13075 8497
rect 11915 8307 11949 8435
rect 13125 8307 13159 8435
rect 11999 8245 13075 8279
rect 10553 8199 11629 8233
rect 10469 8003 10503 8171
rect 11679 8003 11713 8171
rect 10553 7941 11629 7975
rect 11999 8103 13075 8137
rect 11915 7947 11949 8075
rect 13125 7947 13159 8075
rect 11999 7885 13075 7919
rect 10553 7775 11629 7809
rect 10469 7579 10503 7747
rect 11679 7579 11713 7747
rect 10553 7517 11629 7551
rect 11999 7743 13075 7777
rect 11915 7587 11949 7715
rect 13125 7587 13159 7715
rect 11999 7525 13075 7559
rect 15117 17732 15155 17766
rect 15055 15977 15089 17673
rect 15183 15977 15217 17673
rect 15117 15884 15155 15918
rect 15534 17386 15635 17554
rect 16250 17462 17426 17496
rect 16166 17288 16200 17434
rect 17476 17288 17510 17434
rect 16250 17226 17426 17260
rect 16250 17092 17426 17126
rect 16166 16918 16200 17064
rect 17476 16918 17510 17064
rect 16250 16856 17426 16890
rect 16548 16694 17136 16728
rect 16486 16324 16520 16644
rect 17164 16324 17198 16644
rect 17436 16622 17614 16656
rect 17374 16432 17408 16572
rect 17642 16432 17676 16572
rect 17436 16348 17614 16382
rect 16548 16240 17136 16274
rect 14994 13468 15148 13502
rect 15494 13468 15648 13502
rect 15994 13468 16148 13502
rect 16494 13468 16648 13502
rect 16994 13468 17148 13502
rect 17494 13468 17648 13502
rect 14901 12694 14935 13440
rect 15207 12694 15241 13440
rect 15401 12694 15435 13440
rect 15707 12694 15741 13440
rect 15901 12694 15935 13440
rect 16207 12694 16241 13440
rect 16401 12694 16435 13440
rect 16707 12694 16741 13440
rect 16901 12694 16935 13440
rect 17207 12694 17241 13440
rect 17401 12694 17435 13440
rect 17707 12694 17741 13440
rect 14994 12632 15148 12666
rect 15494 12632 15648 12666
rect 15994 12632 16148 12666
rect 16494 12632 16648 12666
rect 16994 12632 17148 12666
rect 17494 12632 17648 12666
rect 18062 12101 18236 13538
rect 14564 11712 14818 11746
rect 14502 10648 14536 11662
rect 14846 10648 14880 11662
rect 14564 10564 14818 10598
rect 14564 10456 14818 10490
rect 14502 9392 14536 10406
rect 14846 9392 14880 10406
rect 14564 9308 14818 9342
rect 17098 11313 18108 11347
rect 17005 11243 17039 11285
rect 18167 11243 18201 11285
rect 17098 11181 18108 11215
rect 17513 10441 17670 10602
rect 17513 10407 17670 10441
rect 17513 10323 17670 10407
rect 17041 10246 18231 10280
rect 16948 9996 16982 10218
rect 18290 9996 18324 10218
rect 17041 9934 18231 9968
rect 17041 9646 18231 9680
rect 16948 9396 16982 9618
rect 18290 9396 18324 9618
rect 17041 9334 18231 9368
rect 14538 8636 14638 8670
rect 14938 8636 15038 8670
rect 15338 8636 15438 8670
rect 15738 8636 15838 8670
rect 16138 8636 16238 8670
rect 16538 8636 16638 8670
rect 16938 8636 17038 8670
rect 17338 8636 17438 8670
rect 17738 8636 17838 8670
rect 18138 8636 18238 8670
rect 14476 7590 14510 8586
rect 14666 7590 14700 8586
rect 14876 7590 14910 8586
rect 15066 7590 15100 8586
rect 15276 7590 15310 8586
rect 15466 7590 15500 8586
rect 15676 7590 15710 8586
rect 15866 7590 15900 8586
rect 16076 7590 16110 8586
rect 16266 7590 16300 8586
rect 16476 7590 16510 8586
rect 16666 7590 16700 8586
rect 16876 7590 16910 8586
rect 17066 7590 17100 8586
rect 17276 7590 17310 8586
rect 17466 7590 17500 8586
rect 17676 7590 17710 8586
rect 17866 7590 17900 8586
rect 18076 7590 18110 8586
rect 18266 7590 18300 8586
rect 14538 7506 14638 7540
rect 14938 7506 15038 7540
rect 15338 7506 15438 7540
rect 15738 7506 15838 7540
rect 16138 7506 16238 7540
rect 16538 7506 16638 7540
rect 16938 7506 17038 7540
rect 17338 7506 17438 7540
rect 17738 7506 17838 7540
rect 18138 7506 18238 7540
<< metal1 >>
rect 6985 19644 10381 19680
rect 6985 19508 7113 19644
rect 10289 19508 10381 19644
rect 6985 19503 10381 19508
rect 1199 19483 2620 19490
rect 1198 19425 2620 19483
rect -81 19029 419 19035
rect -81 18995 -69 19029
rect 407 18995 419 19029
rect -81 18989 419 18995
rect -159 18967 -113 18979
rect -159 18799 -153 18967
rect -119 18799 -113 18967
rect -159 18783 -113 18799
rect 451 18967 497 18979
rect 451 18799 457 18967
rect 491 18799 497 18967
rect 451 18787 497 18799
rect -81 18771 419 18777
rect -81 18737 -69 18771
rect 407 18737 419 18771
rect 1198 18753 1251 19425
rect 1390 19279 1782 19285
rect 1390 19245 1402 19279
rect 1770 19245 1782 19279
rect 1390 19239 1782 19245
rect 2090 19279 2482 19285
rect 2090 19245 2102 19279
rect 2470 19245 2482 19279
rect 2090 19239 2482 19245
rect 1334 19186 1380 19198
rect 1334 19110 1340 19186
rect 1374 19110 1380 19186
rect 1334 19098 1380 19110
rect 1792 19186 1838 19198
rect 1792 19110 1798 19186
rect 1832 19110 1838 19186
rect 1792 19098 1838 19110
rect 2034 19186 2080 19198
rect 2034 19110 2040 19186
rect 2074 19110 2080 19186
rect 2034 19098 2080 19110
rect 2492 19186 2538 19198
rect 2492 19110 2498 19186
rect 2532 19110 2538 19186
rect 2492 19098 2538 19110
rect 1390 19051 1782 19057
rect 1390 19017 1402 19051
rect 1770 19017 1782 19051
rect 1390 19011 1782 19017
rect 2090 19051 2482 19057
rect 2090 19017 2102 19051
rect 2470 19017 2482 19051
rect 2090 19011 2482 19017
rect 2588 18901 2620 19425
rect 5797 19470 11839 19503
rect 3086 19295 3478 19301
rect 3086 19261 3098 19295
rect 3466 19261 3478 19295
rect 3086 19255 3478 19261
rect 3786 19295 4178 19301
rect 3786 19261 3798 19295
rect 4166 19261 4178 19295
rect 3786 19255 4178 19261
rect 5797 19267 5839 19470
rect 5895 19339 6047 19345
rect 5895 19305 5907 19339
rect 6035 19305 6047 19339
rect 5895 19299 6047 19305
rect 6197 19267 6239 19470
rect 6295 19339 6447 19345
rect 6295 19305 6307 19339
rect 6435 19305 6447 19339
rect 6295 19299 6447 19305
rect 6597 19267 6639 19470
rect 6695 19339 6847 19345
rect 6695 19305 6707 19339
rect 6835 19305 6847 19339
rect 6695 19299 6847 19305
rect 6997 19267 7039 19470
rect 7095 19339 7247 19345
rect 7095 19305 7107 19339
rect 7235 19305 7247 19339
rect 7095 19299 7247 19305
rect 7397 19267 7439 19470
rect 7495 19339 7647 19345
rect 7495 19305 7507 19339
rect 7635 19305 7647 19339
rect 7495 19299 7647 19305
rect 7797 19267 7839 19470
rect 7895 19339 8047 19345
rect 7895 19305 7907 19339
rect 8035 19305 8047 19339
rect 7895 19299 8047 19305
rect 8197 19267 8239 19470
rect 8295 19339 8447 19345
rect 8295 19305 8307 19339
rect 8435 19305 8447 19339
rect 8295 19299 8447 19305
rect 8597 19267 8639 19470
rect 8695 19339 8847 19345
rect 8695 19305 8707 19339
rect 8835 19305 8847 19339
rect 8695 19299 8847 19305
rect 8997 19267 9039 19470
rect 9095 19339 9247 19345
rect 9095 19305 9107 19339
rect 9235 19305 9247 19339
rect 9095 19299 9247 19305
rect 9397 19267 9439 19470
rect 9495 19339 9647 19345
rect 9495 19305 9507 19339
rect 9635 19305 9647 19339
rect 9495 19299 9647 19305
rect 9797 19267 9839 19470
rect 9895 19339 10047 19345
rect 9895 19305 9907 19339
rect 10035 19305 10047 19339
rect 9895 19299 10047 19305
rect 10197 19267 10239 19470
rect 10295 19339 10447 19345
rect 10295 19305 10307 19339
rect 10435 19305 10447 19339
rect 10295 19299 10447 19305
rect 10597 19267 10639 19470
rect 10695 19339 10847 19345
rect 10695 19305 10707 19339
rect 10835 19305 10847 19339
rect 10695 19299 10847 19305
rect 10997 19267 11039 19470
rect 11095 19339 11247 19345
rect 11095 19305 11107 19339
rect 11235 19305 11247 19339
rect 11095 19299 11247 19305
rect 11397 19267 11439 19470
rect 11495 19339 11647 19345
rect 11495 19305 11507 19339
rect 11635 19305 11647 19339
rect 11495 19299 11647 19305
rect 11797 19267 11839 19470
rect 11895 19339 12047 19345
rect 11895 19305 11907 19339
rect 12035 19305 12047 19339
rect 11895 19299 12047 19305
rect 5797 19255 5885 19267
rect 3030 19202 3076 19214
rect 3030 19126 3036 19202
rect 3070 19126 3076 19202
rect 3030 19114 3076 19126
rect 3488 19202 3534 19214
rect 3488 19126 3494 19202
rect 3528 19126 3534 19202
rect 3488 19114 3534 19126
rect 3730 19202 3776 19214
rect 3730 19126 3736 19202
rect 3770 19126 3776 19202
rect 3730 19114 3776 19126
rect 4188 19202 4234 19214
rect 4188 19126 4194 19202
rect 4228 19126 4234 19202
rect 4188 19114 4234 19126
rect 3086 19067 3478 19073
rect 3086 19033 3098 19067
rect 3466 19033 3478 19067
rect 3086 19027 3478 19033
rect 3786 19067 4178 19073
rect 3786 19033 3798 19067
rect 4166 19033 4178 19067
rect 3786 19027 4178 19033
rect 1390 18895 1782 18901
rect 1390 18861 1402 18895
rect 1770 18861 1782 18895
rect 1390 18855 1782 18861
rect 2090 18895 2620 18901
rect 2090 18861 2102 18895
rect 2470 18861 2620 18895
rect 2090 18855 2620 18861
rect -81 18731 419 18737
rect 1137 18718 1251 18753
rect -332 18622 419 18654
rect -333 18613 419 18622
rect -333 18601 -69 18613
rect -333 15580 -267 18601
rect -81 18579 -69 18601
rect 407 18579 419 18613
rect -81 18573 419 18579
rect -159 18551 -113 18567
rect -159 18383 -153 18551
rect -119 18383 -113 18551
rect -159 18135 -113 18383
rect 451 18551 497 18563
rect 451 18383 457 18551
rect 491 18383 497 18551
rect 1137 18558 1151 18718
rect 1234 18633 1251 18718
rect 1334 18802 1380 18814
rect 1334 18633 1340 18802
rect 1234 18558 1340 18633
rect 1137 18527 1340 18558
rect 1200 18526 1340 18527
rect 451 18371 497 18383
rect -81 18355 419 18361
rect -81 18321 -69 18355
rect 407 18321 419 18355
rect -81 18315 419 18321
rect 1334 18326 1340 18526
rect 1374 18326 1380 18802
rect 1334 18314 1380 18326
rect 1792 18802 1838 18814
rect 1792 18326 1798 18802
rect 1832 18624 1838 18802
rect 2034 18802 2080 18814
rect 2034 18624 2040 18802
rect 1832 18603 2040 18624
rect 1832 18539 1898 18603
rect 1954 18539 2040 18603
rect 1832 18517 2040 18539
rect 1832 18326 1838 18517
rect 1792 18314 1838 18326
rect 1390 18267 1782 18273
rect -81 18199 837 18249
rect -81 18197 419 18199
rect -81 18163 -69 18197
rect 407 18163 419 18197
rect -81 18157 419 18163
rect -159 17967 -153 18135
rect -119 17967 -113 18135
rect -159 17719 -113 17967
rect 451 18135 497 18147
rect 451 17967 457 18135
rect 491 17967 497 18135
rect 451 17955 497 17967
rect -81 17939 419 17945
rect -81 17905 -69 17939
rect 407 17905 419 17939
rect -81 17899 419 17905
rect -81 17783 543 17833
rect -81 17781 419 17783
rect -81 17747 -69 17781
rect 407 17747 419 17781
rect -81 17741 419 17747
rect 497 17731 543 17783
rect -159 17551 -153 17719
rect -119 17551 -113 17719
rect -159 17303 -113 17551
rect 451 17719 543 17731
rect 451 17551 457 17719
rect 491 17674 543 17719
rect 491 17606 680 17674
rect 491 17551 548 17606
rect 451 17539 548 17551
rect -81 17523 419 17529
rect -81 17489 -69 17523
rect 407 17489 419 17523
rect -81 17483 419 17489
rect 497 17417 548 17539
rect -81 17367 548 17417
rect -81 17365 419 17367
rect -81 17331 -69 17365
rect 407 17331 419 17365
rect -81 17325 419 17331
rect 497 17358 548 17367
rect 649 17358 680 17606
rect 497 17315 680 17358
rect -159 17135 -153 17303
rect -119 17135 -113 17303
rect -159 16887 -113 17135
rect 451 17303 680 17315
rect 451 17135 457 17303
rect 491 17298 680 17303
rect 764 17473 837 18199
rect 1390 18233 1402 18267
rect 1770 18233 1782 18267
rect 1390 18111 1782 18233
rect 1390 18077 1402 18111
rect 1770 18077 1782 18111
rect 1390 18071 1782 18077
rect 1274 18018 1380 18030
rect 1274 17542 1340 18018
rect 1374 17542 1380 18018
rect 1274 17530 1380 17542
rect 1792 18018 1838 18030
rect 1792 17542 1798 18018
rect 1832 17542 1838 18018
rect 1792 17530 1838 17542
rect 1274 17473 1334 17530
rect 764 17326 1334 17473
rect 491 17135 543 17298
rect 451 17123 543 17135
rect -81 17107 419 17113
rect -81 17073 -69 17107
rect 407 17073 419 17107
rect -81 17067 419 17073
rect 764 17001 837 17326
rect -81 16951 837 17001
rect -81 16949 419 16951
rect -81 16915 -69 16949
rect 407 16915 419 16949
rect -81 16909 419 16915
rect -159 16719 -153 16887
rect -119 16719 -113 16887
rect -159 16471 -113 16719
rect 451 16887 497 16899
rect 451 16719 457 16887
rect 491 16719 497 16887
rect 451 16707 497 16719
rect -81 16691 419 16697
rect -81 16657 -69 16691
rect 407 16657 419 16691
rect -81 16651 419 16657
rect 618 16585 681 16587
rect -81 16535 681 16585
rect -81 16533 419 16535
rect -81 16499 -69 16533
rect 407 16499 419 16533
rect -81 16493 419 16499
rect -159 16303 -153 16471
rect -119 16303 -113 16471
rect -159 16287 -113 16303
rect 451 16471 497 16483
rect 451 16303 457 16471
rect 491 16303 497 16471
rect 451 16291 497 16303
rect -81 16275 419 16281
rect -81 16241 -69 16275
rect 407 16241 419 16275
rect -81 16235 419 16241
rect -81 16117 419 16123
rect -81 16083 -69 16117
rect 407 16083 419 16117
rect -81 16077 419 16083
rect -159 16055 -113 16071
rect -159 15887 -153 16055
rect -119 15887 -113 16055
rect -159 15875 -113 15887
rect 451 16055 497 16067
rect 451 15887 457 16055
rect 491 15887 497 16055
rect 451 15875 497 15887
rect -81 15859 419 15865
rect -81 15825 -69 15859
rect 407 15825 419 15859
rect -81 15819 419 15825
rect -345 15575 -23 15580
rect 618 15575 681 16535
rect -345 15546 681 15575
rect -345 15349 -320 15546
rect -55 15476 681 15546
rect -55 15349 -23 15476
rect 769 15367 837 16951
rect 1274 17246 1334 17326
rect 1390 17483 1782 17489
rect 1390 17449 1402 17483
rect 1770 17449 1782 17483
rect 1390 17327 1782 17449
rect 1390 17293 1402 17327
rect 1770 17293 1782 17327
rect 1390 17287 1782 17293
rect 1274 17234 1380 17246
rect 1274 16758 1340 17234
rect 1374 16758 1380 17234
rect 1274 16746 1380 16758
rect 1792 17234 1838 17246
rect 1792 16758 1798 17234
rect 1832 16758 1838 17234
rect 1792 16746 1838 16758
rect 1390 16699 1782 16705
rect 1390 16665 1402 16699
rect 1770 16665 1782 16699
rect 1390 16543 1782 16665
rect 1390 16509 1402 16543
rect 1770 16509 1782 16543
rect 1390 16503 1782 16509
rect 1334 16450 1380 16462
rect 1135 16351 1249 16384
rect 1135 16308 1148 16351
rect -345 15320 -23 15349
rect 149 15281 837 15367
rect 922 16197 1148 16308
rect 149 14992 215 15281
rect 922 15071 1016 16197
rect 1135 16191 1148 16197
rect 1231 16266 1249 16351
rect 1334 16267 1340 16450
rect 1282 16266 1340 16267
rect 1231 16191 1340 16266
rect 1135 16160 1340 16191
rect 1135 16158 1249 16160
rect 1334 15974 1340 16160
rect 1374 15974 1380 16450
rect 1149 15945 1278 15964
rect 1334 15962 1380 15974
rect 1792 16450 1838 16462
rect 1792 15974 1798 16450
rect 1832 16263 1838 16450
rect 1887 16263 1965 18517
rect 2034 18326 2040 18517
rect 2074 18326 2080 18802
rect 2034 18314 2080 18326
rect 2492 18802 2538 18814
rect 2492 18326 2498 18802
rect 2532 18326 2538 18802
rect 2492 18314 2538 18326
rect 2588 18273 2620 18855
rect 2090 18267 2620 18273
rect 2090 18233 2102 18267
rect 2470 18233 2620 18267
rect 2090 18227 2620 18233
rect 2588 18117 2620 18227
rect 2090 18111 2620 18117
rect 2090 18077 2102 18111
rect 2470 18077 2620 18111
rect 2090 18071 2620 18077
rect 2034 18018 2080 18030
rect 2034 17542 2040 18018
rect 2074 17542 2080 18018
rect 2034 17530 2080 17542
rect 2492 18018 2538 18030
rect 2492 17542 2498 18018
rect 2532 17542 2538 18018
rect 2492 17530 2538 17542
rect 2588 17489 2620 18071
rect 2090 17483 2620 17489
rect 2090 17449 2102 17483
rect 2470 17449 2620 17483
rect 2090 17443 2620 17449
rect 2588 17333 2620 17443
rect 2090 17327 2620 17333
rect 2090 17293 2102 17327
rect 2470 17293 2620 17327
rect 2090 17287 2620 17293
rect 2034 17234 2080 17246
rect 2034 16758 2040 17234
rect 2074 16758 2080 17234
rect 2034 16746 2080 16758
rect 2492 17234 2538 17246
rect 2492 16758 2498 17234
rect 2532 16758 2538 17234
rect 2492 16746 2538 16758
rect 2588 16705 2620 17287
rect 2090 16699 2620 16705
rect 2090 16665 2102 16699
rect 2470 16665 2620 16699
rect 2090 16659 2620 16665
rect 2588 16549 2620 16659
rect 2090 16543 2620 16549
rect 2090 16509 2102 16543
rect 2470 16509 2620 16543
rect 2090 16503 2620 16509
rect 2034 16450 2080 16462
rect 2034 16263 2040 16450
rect 1832 16241 2040 16263
rect 1832 16177 1901 16241
rect 1957 16177 2040 16241
rect 1832 16156 2040 16177
rect 1832 15974 1838 16156
rect 1792 15962 1838 15974
rect 2034 15974 2040 16156
rect 2074 15974 2080 16450
rect 2034 15962 2080 15974
rect 2492 16450 2538 16462
rect 2492 15974 2498 16450
rect 2532 15974 2538 16450
rect 2492 15962 2538 15974
rect 1149 15765 1167 15945
rect 1256 15765 1278 15945
rect 2588 15921 2620 16503
rect 1390 15915 1782 15921
rect 1390 15881 1402 15915
rect 1770 15881 1782 15915
rect 1390 15875 1782 15881
rect 2090 15915 2620 15921
rect 2090 15881 2102 15915
rect 2470 15881 2620 15915
rect 2090 15875 2620 15881
rect 2747 18911 3479 18955
rect 2747 18895 3098 18911
rect 1149 15735 1278 15765
rect 1390 15759 1782 15765
rect 1173 15332 1243 15735
rect 1390 15725 1402 15759
rect 1770 15725 1782 15759
rect 1390 15719 1782 15725
rect 2090 15759 2482 15765
rect 2090 15725 2102 15759
rect 2470 15725 2482 15759
rect 2090 15719 2482 15725
rect 1334 15666 1380 15678
rect 1334 15590 1340 15666
rect 1374 15590 1380 15666
rect 1334 15578 1380 15590
rect 1792 15666 1838 15678
rect 1792 15590 1798 15666
rect 1832 15590 1838 15666
rect 1792 15578 1838 15590
rect 2034 15666 2080 15678
rect 2034 15590 2040 15666
rect 2074 15590 2080 15666
rect 2034 15578 2080 15590
rect 2492 15666 2538 15678
rect 2492 15590 2498 15666
rect 2532 15590 2538 15666
rect 2492 15578 2538 15590
rect 1390 15531 1782 15537
rect 1390 15497 1402 15531
rect 1770 15497 1782 15531
rect 1390 15491 1782 15497
rect 2090 15531 2482 15537
rect 2090 15497 2102 15531
rect 2470 15497 2482 15531
rect 2090 15491 2482 15497
rect 2747 15332 2815 18895
rect 3086 18877 3098 18895
rect 3466 18895 3479 18911
rect 3786 18911 4178 18917
rect 3466 18877 3478 18895
rect 3086 18871 3478 18877
rect 3786 18877 3798 18911
rect 4166 18877 4178 18911
rect 3786 18871 4178 18877
rect 2987 18818 3076 18830
rect 2987 18342 3036 18818
rect 3070 18342 3076 18818
rect 2987 18330 3076 18342
rect 3488 18818 3534 18830
rect 3488 18342 3494 18818
rect 3528 18646 3534 18818
rect 3730 18818 3776 18830
rect 3730 18646 3736 18818
rect 3528 18519 3736 18646
rect 3528 18342 3534 18519
rect 3488 18330 3534 18342
rect 2987 18046 3030 18330
rect 3086 18283 3478 18289
rect 3086 18249 3098 18283
rect 3466 18249 3478 18283
rect 3086 18127 3478 18249
rect 3086 18093 3098 18127
rect 3466 18093 3478 18127
rect 3086 18087 3478 18093
rect 2934 18034 3076 18046
rect 2934 17963 3036 18034
rect 2934 16051 2954 17963
rect 3006 17558 3036 17963
rect 3070 17558 3076 18034
rect 3006 17546 3076 17558
rect 3488 18034 3534 18046
rect 3488 17558 3494 18034
rect 3528 17862 3534 18034
rect 3593 17862 3658 18519
rect 3730 18342 3736 18519
rect 3770 18342 3776 18818
rect 3730 18330 3776 18342
rect 4188 18818 4234 18830
rect 4188 18342 4194 18818
rect 4228 18342 4234 18818
rect 4188 18330 4234 18342
rect 3786 18283 4178 18289
rect 3786 18249 3798 18283
rect 4166 18249 4178 18283
rect 3786 18127 4178 18249
rect 5797 18179 5845 19255
rect 5879 18179 5885 19255
rect 5797 18167 5885 18179
rect 6057 19255 6145 19267
rect 6057 18179 6063 19255
rect 6097 18179 6145 19255
rect 6057 18167 6145 18179
rect 6197 19255 6285 19267
rect 6197 18179 6245 19255
rect 6279 18179 6285 19255
rect 6197 18167 6285 18179
rect 6457 19255 6545 19267
rect 6457 18179 6463 19255
rect 6497 18179 6545 19255
rect 6457 18167 6545 18179
rect 6597 19255 6685 19267
rect 6597 18179 6645 19255
rect 6679 18179 6685 19255
rect 6597 18167 6685 18179
rect 6857 19255 6945 19267
rect 6857 18179 6863 19255
rect 6897 18179 6945 19255
rect 6857 18167 6945 18179
rect 6997 19255 7085 19267
rect 6997 18179 7045 19255
rect 7079 18179 7085 19255
rect 6997 18167 7085 18179
rect 7257 19255 7345 19267
rect 7257 18179 7263 19255
rect 7297 18179 7345 19255
rect 7257 18167 7345 18179
rect 7397 19255 7485 19267
rect 7397 18179 7445 19255
rect 7479 18179 7485 19255
rect 7397 18167 7485 18179
rect 7657 19255 7745 19267
rect 7657 18179 7663 19255
rect 7697 18179 7745 19255
rect 7657 18167 7745 18179
rect 7797 19255 7885 19267
rect 7797 18179 7845 19255
rect 7879 18179 7885 19255
rect 7797 18167 7885 18179
rect 8057 19255 8145 19267
rect 8057 18179 8063 19255
rect 8097 18179 8145 19255
rect 8057 18167 8145 18179
rect 8197 19255 8285 19267
rect 8197 18179 8245 19255
rect 8279 18179 8285 19255
rect 8197 18167 8285 18179
rect 8457 19255 8545 19267
rect 8457 18179 8463 19255
rect 8497 18179 8545 19255
rect 8457 18167 8545 18179
rect 8597 19255 8685 19267
rect 8597 18179 8645 19255
rect 8679 18179 8685 19255
rect 8597 18167 8685 18179
rect 8857 19255 8945 19267
rect 8857 18179 8863 19255
rect 8897 18179 8945 19255
rect 8857 18167 8945 18179
rect 8997 19255 9085 19267
rect 8997 18179 9045 19255
rect 9079 18179 9085 19255
rect 8997 18167 9085 18179
rect 9257 19255 9345 19267
rect 9257 18179 9263 19255
rect 9297 18179 9345 19255
rect 9257 18167 9345 18179
rect 9397 19255 9485 19267
rect 9397 18179 9445 19255
rect 9479 18179 9485 19255
rect 9397 18167 9485 18179
rect 9657 19255 9745 19267
rect 9657 18179 9663 19255
rect 9697 18179 9745 19255
rect 9657 18167 9745 18179
rect 9797 19255 9885 19267
rect 9797 18179 9845 19255
rect 9879 18179 9885 19255
rect 9797 18167 9885 18179
rect 10057 19255 10145 19267
rect 10057 18179 10063 19255
rect 10097 18179 10145 19255
rect 10057 18167 10145 18179
rect 10197 19255 10285 19267
rect 10197 18179 10245 19255
rect 10279 18179 10285 19255
rect 10197 18167 10285 18179
rect 10457 19255 10545 19267
rect 10457 18179 10463 19255
rect 10497 18179 10545 19255
rect 10457 18167 10545 18179
rect 10597 19255 10685 19267
rect 10597 18179 10645 19255
rect 10679 18179 10685 19255
rect 10597 18167 10685 18179
rect 10857 19255 10945 19267
rect 10857 18179 10863 19255
rect 10897 18179 10945 19255
rect 10857 18167 10945 18179
rect 10997 19255 11085 19267
rect 10997 18179 11045 19255
rect 11079 18179 11085 19255
rect 10997 18167 11085 18179
rect 11257 19255 11345 19267
rect 11257 18179 11263 19255
rect 11297 18179 11345 19255
rect 11257 18167 11345 18179
rect 11397 19255 11485 19267
rect 11397 18179 11445 19255
rect 11479 18179 11485 19255
rect 11397 18167 11485 18179
rect 11657 19255 11745 19267
rect 11657 18179 11663 19255
rect 11697 18179 11745 19255
rect 11657 18167 11745 18179
rect 11797 19255 11885 19267
rect 11797 18179 11845 19255
rect 11879 18179 11885 19255
rect 11797 18167 11885 18179
rect 12057 19255 12145 19267
rect 12057 18179 12063 19255
rect 12097 18179 12145 19255
rect 12057 18167 12145 18179
rect 3786 18093 3798 18127
rect 4166 18093 4178 18127
rect 3786 18087 4178 18093
rect 5895 18129 6047 18135
rect 5895 18095 5907 18129
rect 6035 18095 6047 18129
rect 5895 18089 6047 18095
rect 3730 18034 3776 18046
rect 3730 17862 3736 18034
rect 3528 17735 3736 17862
rect 3528 17558 3534 17735
rect 3488 17546 3534 17558
rect 3006 17262 3030 17546
rect 3086 17499 3478 17505
rect 3086 17465 3098 17499
rect 3466 17465 3478 17499
rect 3086 17343 3478 17465
rect 3086 17309 3098 17343
rect 3466 17309 3478 17343
rect 3086 17303 3478 17309
rect 3006 17250 3076 17262
rect 3006 16774 3036 17250
rect 3070 16774 3076 17250
rect 3006 16762 3076 16774
rect 3488 17250 3534 17262
rect 3488 16774 3494 17250
rect 3528 17078 3534 17250
rect 3593 17078 3658 17735
rect 3730 17558 3736 17735
rect 3770 17558 3776 18034
rect 3730 17546 3776 17558
rect 4188 18034 4234 18046
rect 4188 17558 4194 18034
rect 4228 17558 4234 18034
rect 6103 17995 6145 18167
rect 6295 18129 6447 18135
rect 6295 18095 6307 18129
rect 6435 18095 6447 18129
rect 6295 18089 6447 18095
rect 6503 17995 6545 18167
rect 6695 18129 6847 18135
rect 6695 18095 6707 18129
rect 6835 18095 6847 18129
rect 6695 18089 6847 18095
rect 6903 17995 6945 18167
rect 7095 18129 7247 18135
rect 7095 18095 7107 18129
rect 7235 18095 7247 18129
rect 7095 18089 7247 18095
rect 7303 17995 7345 18167
rect 7495 18129 7647 18135
rect 7495 18095 7507 18129
rect 7635 18095 7647 18129
rect 7495 18089 7647 18095
rect 7703 17995 7745 18167
rect 7895 18129 8047 18135
rect 7895 18095 7907 18129
rect 8035 18095 8047 18129
rect 7895 18089 8047 18095
rect 8103 17995 8145 18167
rect 8295 18129 8447 18135
rect 8295 18095 8307 18129
rect 8435 18095 8447 18129
rect 8295 18089 8447 18095
rect 8503 17995 8545 18167
rect 8695 18129 8847 18135
rect 8695 18095 8707 18129
rect 8835 18095 8847 18129
rect 8695 18089 8847 18095
rect 8903 17995 8945 18167
rect 9095 18129 9247 18135
rect 9095 18095 9107 18129
rect 9235 18095 9247 18129
rect 9095 18089 9247 18095
rect 9303 17995 9345 18167
rect 9495 18129 9647 18135
rect 9495 18095 9507 18129
rect 9635 18095 9647 18129
rect 9495 18089 9647 18095
rect 9703 17995 9745 18167
rect 9895 18129 10047 18135
rect 9895 18095 9907 18129
rect 10035 18095 10047 18129
rect 9895 18089 10047 18095
rect 10103 17995 10145 18167
rect 10295 18129 10447 18135
rect 10295 18095 10307 18129
rect 10435 18095 10447 18129
rect 10295 18089 10447 18095
rect 10503 17995 10545 18167
rect 10695 18129 10847 18135
rect 10695 18095 10707 18129
rect 10835 18095 10847 18129
rect 10695 18089 10847 18095
rect 10903 17995 10945 18167
rect 11095 18129 11247 18135
rect 11095 18095 11107 18129
rect 11235 18095 11247 18129
rect 11095 18089 11247 18095
rect 11303 17995 11345 18167
rect 11495 18129 11647 18135
rect 11495 18095 11507 18129
rect 11635 18095 11647 18129
rect 11495 18089 11647 18095
rect 11703 17995 11745 18167
rect 11895 18129 12047 18135
rect 11895 18095 11907 18129
rect 12035 18095 12047 18129
rect 11895 18089 12047 18095
rect 12103 17995 12145 18167
rect 6103 17992 12145 17995
rect 6103 17962 12417 17992
rect 11103 17945 12417 17962
rect 10069 17815 10561 17846
rect 10069 17805 10110 17815
rect 9734 17804 10110 17805
rect 7840 17803 10110 17804
rect 4188 17546 4234 17558
rect 5676 17774 10110 17803
rect 5676 17770 8518 17774
rect 5676 17567 5718 17770
rect 5774 17639 5926 17645
rect 5774 17605 5786 17639
rect 5914 17605 5926 17639
rect 5774 17599 5926 17605
rect 6076 17567 6118 17770
rect 6174 17639 6326 17645
rect 6174 17605 6186 17639
rect 6314 17605 6326 17639
rect 6174 17599 6326 17605
rect 6476 17567 6518 17770
rect 6574 17639 6726 17645
rect 6574 17605 6586 17639
rect 6714 17605 6726 17639
rect 6574 17599 6726 17605
rect 6876 17567 6918 17770
rect 6974 17639 7126 17645
rect 6974 17605 6986 17639
rect 7114 17605 7126 17639
rect 6974 17599 7126 17605
rect 7276 17567 7318 17770
rect 7374 17639 7526 17645
rect 7374 17605 7386 17639
rect 7514 17605 7526 17639
rect 7374 17599 7526 17605
rect 7676 17567 7718 17770
rect 7774 17639 7926 17645
rect 7774 17605 7786 17639
rect 7914 17605 7926 17639
rect 7774 17599 7926 17605
rect 8076 17567 8118 17770
rect 8174 17639 8326 17645
rect 8174 17605 8186 17639
rect 8314 17605 8326 17639
rect 8174 17599 8326 17605
rect 8476 17567 8518 17770
rect 9635 17734 10110 17774
rect 8574 17639 8726 17645
rect 8574 17605 8586 17639
rect 8714 17605 8726 17639
rect 8574 17599 8726 17605
rect 5676 17555 5764 17567
rect 3786 17499 4178 17505
rect 3786 17465 3798 17499
rect 4166 17465 4178 17499
rect 3786 17343 4178 17465
rect 3786 17309 3798 17343
rect 4166 17309 4178 17343
rect 3786 17303 4178 17309
rect 3730 17250 3776 17262
rect 3730 17078 3736 17250
rect 3528 16951 3736 17078
rect 3528 16774 3534 16951
rect 3488 16762 3534 16774
rect 3006 16478 3030 16762
rect 3086 16715 3478 16721
rect 3086 16681 3098 16715
rect 3466 16681 3478 16715
rect 3086 16559 3478 16681
rect 3086 16525 3098 16559
rect 3466 16525 3478 16559
rect 3086 16519 3478 16525
rect 3006 16466 3076 16478
rect 3006 16051 3036 16466
rect 2934 15990 3036 16051
rect 3070 15990 3076 16466
rect 2934 15978 3076 15990
rect 3488 16466 3534 16478
rect 3488 15990 3494 16466
rect 3528 16294 3534 16466
rect 3593 16294 3658 16951
rect 3730 16774 3736 16951
rect 3770 16774 3776 17250
rect 3730 16762 3776 16774
rect 4188 17250 4234 17262
rect 4188 16774 4194 17250
rect 4228 16774 4234 17250
rect 4188 16762 4234 16774
rect 3786 16715 4178 16721
rect 3786 16681 3798 16715
rect 4166 16681 4178 16715
rect 3786 16559 4178 16681
rect 3786 16525 3798 16559
rect 4166 16525 4178 16559
rect 3786 16519 4178 16525
rect 5676 16479 5724 17555
rect 5758 16479 5764 17555
rect 3730 16466 3776 16478
rect 3730 16294 3736 16466
rect 3528 16167 3736 16294
rect 3528 15990 3534 16167
rect 3488 15978 3534 15990
rect 1173 15264 2815 15332
rect 2987 15694 3030 15978
rect 3086 15931 3478 15937
rect 3086 15897 3098 15931
rect 3466 15897 3478 15931
rect 3086 15775 3478 15897
rect 3086 15741 3098 15775
rect 3466 15741 3478 15775
rect 3086 15735 3478 15741
rect 2987 15682 3076 15694
rect 2987 15206 3036 15682
rect 3070 15206 3076 15682
rect 2987 15194 3076 15206
rect 3488 15682 3534 15694
rect 3488 15206 3494 15682
rect 3528 15510 3534 15682
rect 3593 15673 3658 16167
rect 3730 15990 3736 16167
rect 3770 15990 3776 16466
rect 3730 15978 3776 15990
rect 4188 16466 4234 16478
rect 5676 16467 5764 16479
rect 5936 17555 6024 17567
rect 5936 16479 5942 17555
rect 5976 16479 6024 17555
rect 5936 16467 6024 16479
rect 6076 17555 6164 17567
rect 6076 16479 6124 17555
rect 6158 16479 6164 17555
rect 6076 16467 6164 16479
rect 6336 17555 6424 17567
rect 6336 16479 6342 17555
rect 6376 16479 6424 17555
rect 6336 16467 6424 16479
rect 6476 17555 6564 17567
rect 6476 16479 6524 17555
rect 6558 16479 6564 17555
rect 6476 16467 6564 16479
rect 6736 17555 6824 17567
rect 6736 16479 6742 17555
rect 6776 16479 6824 17555
rect 6736 16467 6824 16479
rect 6876 17555 6964 17567
rect 6876 16479 6924 17555
rect 6958 16479 6964 17555
rect 6876 16467 6964 16479
rect 7136 17555 7224 17567
rect 7136 16479 7142 17555
rect 7176 16479 7224 17555
rect 7136 16467 7224 16479
rect 7276 17555 7364 17567
rect 7276 16479 7324 17555
rect 7358 16479 7364 17555
rect 7276 16467 7364 16479
rect 7536 17555 7624 17567
rect 7536 16479 7542 17555
rect 7576 16479 7624 17555
rect 7536 16467 7624 16479
rect 7676 17555 7764 17567
rect 7676 16479 7724 17555
rect 7758 16479 7764 17555
rect 7676 16467 7764 16479
rect 7936 17555 8024 17567
rect 7936 16479 7942 17555
rect 7976 16479 8024 17555
rect 7936 16467 8024 16479
rect 8076 17555 8164 17567
rect 8076 16479 8124 17555
rect 8158 16479 8164 17555
rect 8076 16467 8164 16479
rect 8336 17555 8424 17567
rect 8336 16479 8342 17555
rect 8376 16479 8424 17555
rect 8336 16467 8424 16479
rect 8476 17555 8564 17567
rect 8476 16479 8524 17555
rect 8558 16479 8564 17555
rect 8476 16467 8564 16479
rect 8736 17555 8824 17567
rect 8736 16479 8742 17555
rect 8776 16479 8824 17555
rect 9635 17522 9761 17734
rect 10069 17718 10110 17734
rect 10525 17718 10561 17815
rect 10069 17698 10561 17718
rect 11103 17720 11162 17945
rect 12344 17720 12417 17945
rect 11103 17676 12417 17720
rect 9314 17482 10074 17522
rect 11819 17490 11935 17676
rect 9314 17314 9362 17482
rect 9418 17395 9570 17401
rect 9418 17361 9430 17395
rect 9558 17361 9570 17395
rect 9418 17355 9570 17361
rect 9818 17395 9970 17401
rect 9818 17361 9830 17395
rect 9958 17361 9970 17395
rect 9818 17355 9970 17361
rect 10026 17314 10074 17482
rect 9314 17302 9408 17314
rect 9314 17126 9368 17302
rect 9402 17126 9408 17302
rect 9314 17114 9408 17126
rect 9580 17302 9626 17314
rect 9580 17126 9586 17302
rect 9620 17126 9626 17302
rect 9580 17114 9626 17126
rect 9762 17302 9808 17314
rect 9762 17126 9768 17302
rect 9802 17126 9808 17302
rect 9762 17114 9808 17126
rect 9980 17302 10074 17314
rect 9980 17126 9986 17302
rect 10020 17161 10074 17302
rect 10579 17452 12127 17490
rect 10579 17285 10621 17452
rect 10677 17366 10829 17372
rect 10677 17332 10689 17366
rect 10817 17332 10829 17366
rect 10677 17326 10829 17332
rect 10979 17285 11021 17452
rect 11077 17366 11229 17372
rect 11077 17332 11089 17366
rect 11217 17332 11229 17366
rect 11077 17326 11229 17332
rect 11477 17366 11629 17372
rect 11477 17332 11489 17366
rect 11617 17332 11629 17366
rect 11477 17326 11629 17332
rect 11685 17285 11727 17452
rect 11877 17366 12029 17372
rect 11877 17332 11889 17366
rect 12017 17332 12029 17366
rect 11877 17326 12029 17332
rect 12085 17285 12127 17452
rect 10579 17273 10667 17285
rect 10020 17126 10186 17161
rect 9980 17114 10186 17126
rect 9418 17067 9970 17073
rect 9418 17033 9430 17067
rect 9558 17033 9830 17067
rect 9958 17033 9970 17067
rect 9418 17027 9970 17033
rect 10121 17045 10186 17114
rect 10579 17097 10627 17273
rect 10661 17097 10667 17273
rect 10579 17085 10667 17097
rect 10839 17273 10935 17285
rect 10839 17097 10845 17273
rect 10879 17097 10935 17273
rect 10839 17085 10935 17097
rect 10979 17273 11067 17285
rect 10979 17097 11027 17273
rect 11061 17097 11067 17273
rect 10979 17085 11067 17097
rect 11239 17273 11285 17285
rect 11239 17097 11245 17273
rect 11279 17144 11285 17273
rect 11421 17273 11467 17285
rect 11421 17144 11427 17273
rect 11279 17097 11427 17144
rect 11461 17097 11467 17273
rect 11239 17085 11467 17097
rect 11639 17273 11727 17285
rect 11639 17097 11645 17273
rect 11679 17097 11727 17273
rect 11639 17085 11727 17097
rect 11771 17273 11867 17285
rect 11771 17097 11827 17273
rect 11861 17097 11867 17273
rect 11771 17085 11867 17097
rect 12039 17273 12127 17285
rect 12039 17097 12045 17273
rect 12079 17097 12127 17273
rect 12039 17085 12127 17097
rect 10121 17044 10711 17045
rect 10121 17038 10829 17044
rect 9457 16628 9520 17027
rect 10121 17004 10689 17038
rect 10817 17004 10829 17038
rect 10121 16998 10829 17004
rect 10885 16890 10935 17085
rect 11077 17038 11229 17044
rect 11077 17004 11089 17038
rect 11217 17004 11229 17038
rect 11077 16998 11229 17004
rect 11328 16890 11378 17085
rect 11477 17038 11629 17044
rect 11477 17004 11489 17038
rect 11617 17004 11629 17038
rect 11477 16998 11629 17004
rect 11771 16890 11821 17085
rect 11877 17038 12029 17044
rect 11877 17004 11889 17038
rect 12017 17004 12029 17038
rect 11877 16998 12029 17004
rect 10885 16851 11821 16890
rect 11150 16762 11180 16851
rect 11520 16762 11543 16851
rect 11150 16748 11543 16762
rect 10509 16692 10811 16723
rect 8736 16467 8824 16479
rect 4188 15990 4194 16466
rect 4228 15990 4234 16466
rect 5774 16429 5926 16435
rect 5774 16395 5786 16429
rect 5914 16395 5926 16429
rect 5774 16389 5926 16395
rect 5982 16295 6024 16467
rect 6174 16429 6326 16435
rect 6174 16395 6186 16429
rect 6314 16395 6326 16429
rect 6174 16389 6326 16395
rect 6382 16295 6424 16467
rect 6574 16429 6726 16435
rect 6574 16395 6586 16429
rect 6714 16395 6726 16429
rect 6574 16389 6726 16395
rect 6782 16295 6824 16467
rect 6974 16429 7126 16435
rect 6974 16395 6986 16429
rect 7114 16395 7126 16429
rect 6974 16389 7126 16395
rect 7182 16295 7224 16467
rect 7374 16429 7526 16435
rect 7374 16395 7386 16429
rect 7514 16395 7526 16429
rect 7374 16389 7526 16395
rect 7582 16295 7624 16467
rect 7774 16429 7926 16435
rect 7774 16395 7786 16429
rect 7914 16395 7926 16429
rect 7774 16389 7926 16395
rect 7982 16295 8024 16467
rect 8174 16429 8326 16435
rect 8174 16395 8186 16429
rect 8314 16395 8326 16429
rect 8174 16389 8326 16395
rect 8382 16295 8424 16467
rect 8574 16429 8726 16435
rect 8574 16395 8586 16429
rect 8714 16395 8726 16429
rect 8574 16389 8726 16395
rect 8782 16295 8824 16467
rect 9010 16574 9850 16628
rect 9010 16473 9084 16574
rect 9010 16375 9052 16473
rect 9786 16379 9850 16574
rect 10509 16388 10546 16692
rect 9594 16375 9850 16379
rect 9010 16343 9850 16375
rect 10508 16377 10546 16388
rect 10771 16388 10811 16692
rect 10771 16377 10812 16388
rect 5982 16264 8824 16295
rect 5982 16262 6477 16264
rect 6419 16165 6477 16262
rect 7983 16262 8824 16264
rect 7983 16165 8021 16262
rect 6419 16143 8021 16165
rect 10508 16088 10812 16377
rect 13052 16088 13638 20761
rect 15556 18292 18647 18571
rect 15055 17766 15217 17782
rect 15055 17732 15117 17766
rect 15155 17732 15217 17766
rect 15105 17726 15167 17732
rect 9473 16082 13638 16088
rect 4188 15978 4234 15990
rect 9336 15974 13638 16082
rect 3786 15931 4178 15937
rect 3786 15897 3798 15931
rect 4166 15897 4178 15931
rect 3786 15775 4178 15897
rect 3786 15741 3798 15775
rect 4166 15741 4178 15775
rect 3786 15735 4178 15741
rect 8388 15724 8672 15725
rect 8388 15707 9189 15724
rect 3593 15510 3598 15673
rect 3528 15391 3598 15510
rect 3653 15510 3658 15673
rect 3730 15682 3776 15694
rect 3730 15510 3736 15682
rect 3653 15391 3736 15510
rect 3528 15383 3736 15391
rect 3528 15206 3534 15383
rect 3488 15194 3534 15206
rect 3730 15206 3736 15383
rect 3770 15206 3776 15682
rect 3730 15194 3776 15206
rect 4188 15682 4234 15694
rect 4188 15206 4194 15682
rect 4228 15206 4234 15682
rect 8388 15638 8416 15707
rect 8643 15638 9189 15707
rect 8388 15635 9189 15638
rect 8388 15625 8672 15635
rect 7125 15561 7330 15603
rect 6450 15527 8801 15561
rect 9130 15558 9189 15635
rect 9336 15598 9383 15974
rect 9629 15851 13638 15974
rect 15049 17673 15095 17685
rect 15049 15977 15055 17673
rect 15089 15977 15095 17673
rect 15049 15965 15095 15977
rect 15177 17673 15223 17685
rect 15177 15977 15183 17673
rect 15217 16381 15223 17673
rect 15556 17580 15835 18292
rect 15505 17554 16508 17580
rect 15505 17386 15534 17554
rect 15635 17502 16508 17554
rect 15635 17500 17438 17502
rect 15635 17386 16060 17500
rect 16238 17496 17438 17500
rect 16238 17462 16250 17496
rect 17426 17462 17438 17496
rect 16238 17456 17438 17462
rect 15505 17362 16060 17386
rect 15914 17174 16060 17362
rect 16104 17434 16206 17446
rect 16104 17288 16114 17434
rect 16200 17288 16206 17434
rect 16104 17276 16206 17288
rect 17470 17434 17660 17446
rect 17470 17288 17476 17434
rect 17562 17288 17660 17434
rect 17470 17276 17660 17288
rect 16238 17260 17438 17266
rect 16238 17226 16250 17260
rect 17426 17226 17438 17260
rect 16238 17220 17438 17226
rect 17382 17214 17438 17220
rect 17572 17214 17590 17276
rect 17382 17178 17590 17214
rect 15914 17132 16508 17174
rect 16238 17126 17438 17132
rect 16238 17092 16250 17126
rect 17426 17092 17438 17126
rect 16238 17086 17438 17092
rect 17572 17078 17590 17178
rect 17646 17078 17660 17276
rect 17572 17076 17660 17078
rect 16104 17064 16206 17076
rect 16104 16918 16114 17064
rect 16200 16918 16206 17064
rect 16104 16906 16206 16918
rect 17470 17064 17660 17076
rect 17470 16918 17476 17064
rect 17562 16918 17660 17064
rect 17470 16906 17660 16918
rect 16104 16780 16146 16906
rect 16238 16890 17438 16896
rect 16238 16856 16250 16890
rect 17426 16856 17438 16890
rect 16238 16850 17438 16856
rect 16238 16780 16346 16850
rect 16104 16732 16346 16780
rect 16238 16570 16346 16732
rect 16536 16804 17148 16850
rect 17584 16804 17660 16906
rect 16536 16754 17660 16804
rect 16536 16728 17148 16754
rect 16536 16694 16548 16728
rect 17136 16694 17148 16728
rect 16536 16688 17148 16694
rect 17424 16656 17660 16754
rect 16480 16644 16526 16656
rect 16480 16570 16486 16644
rect 16238 16406 16486 16570
rect 15770 16381 16016 16396
rect 15217 16370 16016 16381
rect 15217 16308 15770 16370
rect 15970 16308 16016 16370
rect 15217 16303 16016 16308
rect 15217 15977 15223 16303
rect 15770 16278 16016 16303
rect 16238 16234 16368 16406
rect 16480 16324 16486 16406
rect 16520 16324 16526 16644
rect 16480 16312 16526 16324
rect 17158 16644 17204 16656
rect 17158 16324 17164 16644
rect 17198 16584 17204 16644
rect 17424 16622 17436 16656
rect 17614 16622 17660 16656
rect 17424 16616 17660 16622
rect 17198 16572 17414 16584
rect 17198 16562 17374 16572
rect 17198 16438 17234 16562
rect 17336 16438 17374 16562
rect 17198 16432 17374 16438
rect 17408 16432 17414 16572
rect 17198 16420 17414 16432
rect 17636 16572 17682 16584
rect 17636 16432 17642 16572
rect 17676 16432 17682 16572
rect 17636 16420 17682 16432
rect 17198 16324 17204 16420
rect 17158 16312 17204 16324
rect 17424 16382 17626 16388
rect 17424 16348 17436 16382
rect 17614 16348 17626 16382
rect 16536 16274 17148 16280
rect 16536 16240 16548 16274
rect 17136 16240 17148 16274
rect 16536 16234 17148 16240
rect 17424 16234 17626 16348
rect 16238 16176 17626 16234
rect 15177 15965 15223 15977
rect 15055 15918 15217 15924
rect 15055 15884 15117 15918
rect 15155 15884 15217 15918
rect 15055 15878 15217 15884
rect 9629 15598 9683 15851
rect 10345 15724 10629 15725
rect 9336 15566 9683 15598
rect 9828 15707 10629 15724
rect 9828 15638 10374 15707
rect 10601 15638 10629 15707
rect 9828 15635 10629 15638
rect 9828 15558 9887 15635
rect 10345 15625 10629 15635
rect 11687 15561 11892 15603
rect 5930 15525 8801 15527
rect 5930 15521 7030 15525
rect 5930 15487 5942 15521
rect 7018 15487 7030 15521
rect 5930 15481 7030 15487
rect 7280 15521 8801 15525
rect 4188 15194 4234 15206
rect 5810 15459 5898 15471
rect 5810 15331 5858 15459
rect 5892 15331 5898 15459
rect 5810 15319 5898 15331
rect 7062 15459 7150 15471
rect 7062 15331 7068 15459
rect 7102 15331 7150 15459
rect 7062 15319 7150 15331
rect 3086 15147 3478 15153
rect 3086 15113 3098 15147
rect 3466 15113 3478 15147
rect -310 14914 215 14992
rect 711 14996 864 15020
rect 711 14940 749 14996
rect 826 14940 864 14996
rect 922 14971 1593 15071
rect 711 14923 864 14940
rect -310 13994 -254 14914
rect 58 14685 250 14691
rect 58 14651 70 14685
rect 238 14651 250 14685
rect 58 14645 250 14651
rect 474 14685 666 14691
rect 474 14651 486 14685
rect 654 14651 666 14685
rect 474 14645 666 14651
rect 711 14613 761 14923
rect 1127 14914 1593 14971
rect 1856 14996 2009 15020
rect 1856 14940 1894 14996
rect 1971 14940 2009 14996
rect 3086 14991 3478 15113
rect 3086 14957 3098 14991
rect 3466 14957 3478 14991
rect 3086 14951 3478 14957
rect 3786 15147 4178 15153
rect 3786 15113 3798 15147
rect 4166 15113 4178 15147
rect 3786 14991 4178 15113
rect 3786 14957 3798 14991
rect 4166 14957 4178 14991
rect 3786 14951 4178 14957
rect 5810 15111 5852 15319
rect 5930 15303 7030 15309
rect 5930 15269 5942 15303
rect 7018 15269 7030 15303
rect 5930 15263 7030 15269
rect 5930 15161 7030 15167
rect 5930 15127 5942 15161
rect 7018 15127 7030 15161
rect 5930 15121 7030 15127
rect 7108 15111 7150 15319
rect 5810 15099 5898 15111
rect 5810 14971 5858 15099
rect 5892 14971 5898 15099
rect 5810 14959 5898 14971
rect 7062 15099 7150 15111
rect 7062 14971 7068 15099
rect 7102 14971 7150 15099
rect 7280 15427 7328 15521
rect 8733 15492 8801 15521
rect 9063 15552 9263 15558
rect 9063 15518 9075 15552
rect 9251 15518 9263 15552
rect 9063 15512 9263 15518
rect 9754 15552 9954 15558
rect 9754 15518 9766 15552
rect 9942 15518 9954 15552
rect 9754 15512 9954 15518
rect 10216 15527 12567 15561
rect 10216 15525 13087 15527
rect 10216 15521 11737 15525
rect 8976 15492 9022 15502
rect 8733 15490 9022 15492
rect 7406 15477 8506 15483
rect 7406 15443 7418 15477
rect 8494 15443 8506 15477
rect 7406 15437 8506 15443
rect 8733 15432 8982 15490
rect 8733 15431 8801 15432
rect 7280 15415 7374 15427
rect 7280 15367 7334 15415
rect 7368 15367 7374 15415
rect 7280 15355 7374 15367
rect 8538 15415 8632 15427
rect 8538 15367 8544 15415
rect 8578 15367 8632 15415
rect 8538 15355 8632 15367
rect 7280 15265 7328 15355
rect 7406 15339 8506 15345
rect 7406 15305 7418 15339
rect 8494 15305 8506 15339
rect 7406 15299 8506 15305
rect 8584 15265 8632 15355
rect 8976 15362 8982 15432
rect 9016 15362 9022 15490
rect 8976 15350 9022 15362
rect 9304 15490 9350 15502
rect 9304 15362 9310 15490
rect 9344 15362 9350 15490
rect 9304 15350 9350 15362
rect 9667 15490 9713 15502
rect 9667 15362 9673 15490
rect 9707 15362 9713 15490
rect 9667 15350 9713 15362
rect 9995 15492 10041 15502
rect 10216 15492 10284 15521
rect 9995 15490 10284 15492
rect 9995 15362 10001 15490
rect 10035 15432 10284 15490
rect 10511 15477 11611 15483
rect 10511 15443 10523 15477
rect 11599 15443 11611 15477
rect 10511 15437 11611 15443
rect 10035 15362 10041 15432
rect 10216 15431 10284 15432
rect 11689 15427 11737 15521
rect 11987 15521 13087 15525
rect 11987 15487 11999 15521
rect 13075 15487 13087 15521
rect 11987 15481 13087 15487
rect 9995 15350 10041 15362
rect 10385 15415 10479 15427
rect 10385 15367 10439 15415
rect 10473 15367 10479 15415
rect 10385 15355 10479 15367
rect 11643 15415 11737 15427
rect 11643 15367 11649 15415
rect 11683 15367 11737 15415
rect 11643 15355 11737 15367
rect 9063 15334 9263 15340
rect 9063 15300 9075 15334
rect 9251 15300 9263 15334
rect 9063 15294 9263 15300
rect 9754 15334 9954 15340
rect 9754 15300 9766 15334
rect 9942 15300 9954 15334
rect 9754 15294 9954 15300
rect 7280 15221 8632 15265
rect 9143 15239 9187 15294
rect 7280 15129 7328 15221
rect 7406 15179 8506 15185
rect 7406 15145 7418 15179
rect 8494 15145 8506 15179
rect 7406 15139 8506 15145
rect 8584 15129 8632 15221
rect 7280 15117 7374 15129
rect 7280 15069 7334 15117
rect 7368 15069 7374 15117
rect 7280 15057 7374 15069
rect 8538 15117 8632 15129
rect 8538 15069 8544 15117
rect 8578 15069 8632 15117
rect 8538 15057 8632 15069
rect 8730 15194 9187 15239
rect 9249 15246 9436 15264
rect 9249 15194 9274 15246
rect 9372 15194 9436 15246
rect 8730 15162 8802 15194
rect 9249 15179 9436 15194
rect 9581 15246 9768 15264
rect 9581 15194 9645 15246
rect 9743 15194 9768 15246
rect 9830 15239 9874 15294
rect 10385 15265 10433 15355
rect 10511 15339 11611 15345
rect 10511 15305 10523 15339
rect 11599 15305 11611 15339
rect 10511 15299 11611 15305
rect 11689 15265 11737 15355
rect 9830 15194 10287 15239
rect 9581 15179 9768 15194
rect 8730 15079 8748 15162
rect 8783 15079 8802 15162
rect 10215 15162 10287 15194
rect 9063 15144 9263 15150
rect 9063 15110 9075 15144
rect 9251 15110 9263 15144
rect 9063 15104 9263 15110
rect 9754 15144 9954 15150
rect 9754 15110 9766 15144
rect 9942 15110 9954 15144
rect 9754 15104 9954 15110
rect 8730 15063 8802 15079
rect 8976 15082 9022 15094
rect 7406 15041 8506 15047
rect 7406 15007 7418 15041
rect 8494 15012 8506 15041
rect 8494 15007 8749 15012
rect 7406 15001 8749 15007
rect 8249 14971 8749 15001
rect 7062 14959 7150 14971
rect 1856 14923 2009 14940
rect 890 14685 1082 14691
rect 890 14651 902 14685
rect 1070 14651 1082 14685
rect 890 14645 1082 14651
rect 1127 14613 1177 14914
rect 1306 14685 1498 14691
rect 1306 14651 1318 14685
rect 1486 14651 1498 14685
rect 1306 14645 1498 14651
rect 1543 14613 1593 14914
rect 1722 14685 1914 14691
rect 1722 14651 1734 14685
rect 1902 14651 1914 14685
rect 1722 14645 1914 14651
rect 1959 14613 2009 14923
rect 3030 14898 3076 14910
rect 2677 14786 2808 14848
rect 2138 14685 2330 14691
rect 2138 14651 2150 14685
rect 2318 14651 2330 14685
rect 2138 14645 2330 14651
rect 2 14601 48 14613
rect 2 14125 8 14601
rect 42 14125 48 14601
rect 2 14113 48 14125
rect 260 14601 306 14613
rect 260 14125 266 14601
rect 300 14125 306 14601
rect 260 14113 306 14125
rect 418 14601 464 14613
rect 418 14125 424 14601
rect 458 14125 464 14601
rect 418 14113 464 14125
rect 676 14601 761 14613
rect 676 14125 682 14601
rect 716 14347 761 14601
rect 834 14601 880 14613
rect 716 14125 722 14347
rect 676 14113 722 14125
rect 834 14125 840 14601
rect 874 14125 880 14601
rect 834 14113 880 14125
rect 1092 14601 1177 14613
rect 1092 14125 1098 14601
rect 1132 14347 1177 14601
rect 1250 14601 1296 14613
rect 1132 14125 1138 14347
rect 1092 14113 1138 14125
rect 1250 14125 1256 14601
rect 1290 14125 1296 14601
rect 1250 14113 1296 14125
rect 1508 14601 1593 14613
rect 1508 14125 1514 14601
rect 1548 14347 1593 14601
rect 1666 14601 1712 14613
rect 1548 14125 1554 14347
rect 1508 14113 1554 14125
rect 1666 14125 1672 14601
rect 1706 14125 1712 14601
rect 1666 14113 1712 14125
rect 1924 14601 2009 14613
rect 1924 14125 1930 14601
rect 1964 14347 2009 14601
rect 2082 14601 2128 14613
rect 1964 14125 1970 14347
rect 1924 14113 1970 14125
rect 2082 14125 2088 14601
rect 2122 14125 2128 14601
rect 2082 14113 2128 14125
rect 2340 14601 2386 14613
rect 2340 14125 2346 14601
rect 2380 14125 2386 14601
rect 2677 14566 2698 14786
rect 2788 14730 2808 14786
rect 2788 14729 2847 14730
rect 3030 14729 3036 14898
rect 2788 14622 3036 14729
rect 2788 14621 2847 14622
rect 2788 14566 2808 14621
rect 2677 14506 2808 14566
rect 3030 14422 3036 14622
rect 3070 14422 3076 14898
rect 3030 14410 3076 14422
rect 3488 14898 3534 14910
rect 3488 14422 3494 14898
rect 3528 14720 3534 14898
rect 3730 14898 3776 14910
rect 3730 14720 3736 14898
rect 3528 14699 3736 14720
rect 3528 14635 3594 14699
rect 3650 14635 3736 14699
rect 3528 14613 3736 14635
rect 3528 14422 3534 14613
rect 3488 14410 3534 14422
rect 3086 14363 3478 14369
rect 3086 14329 3098 14363
rect 3466 14329 3478 14363
rect 3086 14207 3478 14329
rect 3086 14173 3098 14207
rect 3466 14173 3478 14207
rect 3086 14167 3478 14173
rect 2340 14113 2386 14125
rect 2983 14114 3076 14126
rect 58 14075 254 14081
rect 58 14041 70 14075
rect 238 14041 254 14075
rect 58 14035 254 14041
rect 474 14075 1914 14081
rect 474 14041 486 14075
rect 654 14041 902 14075
rect 1070 14041 1318 14075
rect 1486 14041 1734 14075
rect 1902 14041 1914 14075
rect 474 14035 1914 14041
rect 2134 14075 2330 14081
rect 2134 14041 2150 14075
rect 2318 14041 2330 14075
rect 2134 14035 2330 14041
rect 511 13994 610 14035
rect -310 13944 610 13994
rect 941 13983 1114 13990
rect 941 13946 964 13983
rect 1084 13973 1114 13983
rect 1084 13946 1905 13973
rect 941 13939 1905 13946
rect 987 13937 1905 13939
rect 463 13817 732 13840
rect 245 13807 732 13817
rect 245 13451 495 13807
rect 663 13801 1655 13807
rect 663 13767 675 13801
rect 1643 13767 1655 13801
rect 663 13761 1655 13767
rect 607 13717 653 13729
rect 607 13541 613 13717
rect 647 13541 653 13717
rect 607 13529 653 13541
rect 1665 13717 1711 13729
rect 1665 13541 1671 13717
rect 1705 13626 1711 13717
rect 1865 13626 1905 13937
rect 2983 13655 3036 14114
rect 1705 13584 1905 13626
rect 2024 13638 3036 13655
rect 3070 13638 3076 14114
rect 2024 13626 3076 13638
rect 3488 14114 3534 14126
rect 3488 13638 3494 14114
rect 3528 13638 3534 14114
rect 3488 13626 3534 13638
rect 2024 13608 3030 13626
rect 1705 13541 1711 13584
rect 1665 13529 1711 13541
rect 663 13491 1655 13497
rect 663 13457 675 13491
rect 1643 13457 1655 13491
rect 663 13451 1655 13457
rect 245 13448 730 13451
rect 293 13418 730 13448
rect 293 13160 479 13418
rect 1154 13218 1398 13251
rect 1154 13160 1185 13218
rect 293 13055 1185 13160
rect 1154 13005 1185 13055
rect 1366 13005 1398 13218
rect 2024 13102 2055 13608
rect 2220 13342 3030 13608
rect 3086 13579 3478 13585
rect 3086 13545 3098 13579
rect 3466 13545 3478 13579
rect 3086 13423 3478 13545
rect 3086 13389 3098 13423
rect 3466 13389 3478 13423
rect 3086 13383 3478 13389
rect 2220 13330 3076 13342
rect 2220 13321 3036 13330
rect 2220 13102 2257 13321
rect 2024 13058 2257 13102
rect 1154 12960 1398 13005
rect -248 12916 367 12959
rect -248 12676 -207 12916
rect -163 12726 237 12732
rect -163 12692 -151 12726
rect 225 12692 237 12726
rect -163 12686 237 12692
rect 326 12676 367 12916
rect 2983 12854 3036 13321
rect 3070 12854 3076 13330
rect 2983 12842 3076 12854
rect 3488 13330 3534 13342
rect 3488 12854 3494 13330
rect 3528 12854 3534 13330
rect 3488 12842 3534 12854
rect 3086 12795 3478 12801
rect 3086 12761 3098 12795
rect 3466 12761 3478 12795
rect 473 12726 873 12732
rect 473 12692 485 12726
rect 861 12692 873 12726
rect 473 12686 873 12692
rect 1109 12726 1509 12732
rect 1109 12692 1121 12726
rect 1497 12692 1509 12726
rect 1109 12686 1509 12692
rect 1745 12726 2145 12732
rect 1745 12692 1757 12726
rect 2133 12692 2145 12726
rect 1745 12686 2145 12692
rect -250 12664 -204 12676
rect -250 12596 -244 12664
rect -210 12596 -204 12664
rect -250 12584 -204 12596
rect 278 12664 432 12676
rect 278 12596 284 12664
rect 318 12596 392 12664
rect 426 12596 432 12664
rect 278 12594 432 12596
rect 237 12584 432 12594
rect 914 12664 1068 12676
rect 914 12596 920 12664
rect 954 12596 1028 12664
rect 1062 12596 1068 12664
rect 914 12584 1068 12596
rect 1550 12664 1704 12676
rect 1550 12596 1556 12664
rect 1590 12596 1664 12664
rect 1698 12596 1704 12664
rect 1550 12584 1704 12596
rect 2186 12664 2232 12676
rect 2186 12596 2192 12664
rect 2226 12596 2232 12664
rect 3086 12639 3478 12761
rect 3086 12605 3098 12639
rect 3466 12605 3478 12639
rect 3086 12599 3478 12605
rect 2186 12584 2232 12596
rect 237 12574 371 12584
rect -163 12568 371 12574
rect -163 12534 -151 12568
rect 225 12534 371 12568
rect -163 12528 371 12534
rect 473 12568 873 12574
rect 473 12534 485 12568
rect 861 12534 873 12568
rect 473 12528 873 12534
rect 44 12409 166 12436
rect 44 12308 62 12409
rect 146 12308 166 12409
rect 339 12342 371 12528
rect 639 12342 696 12528
rect 974 12342 1006 12584
rect 1109 12568 1509 12574
rect 1109 12534 1121 12568
rect 1497 12534 1509 12568
rect 1109 12528 1509 12534
rect 1282 12342 1339 12528
rect 1609 12342 1641 12584
rect 1745 12568 2145 12574
rect 1745 12534 1757 12568
rect 2133 12534 2145 12568
rect 1745 12528 2145 12534
rect 1925 12342 1982 12528
rect 2189 12356 2221 12584
rect 3030 12546 3076 12558
rect 2678 12384 2809 12446
rect 2184 12342 2515 12356
rect 44 10997 166 12308
rect 262 12331 2515 12342
rect 262 12273 2207 12331
rect 499 11877 556 12273
rect 2184 12260 2207 12273
rect 2491 12260 2515 12331
rect 2184 12237 2515 12260
rect 2678 12164 2699 12384
rect 2789 12363 2809 12384
rect 3030 12363 3036 12546
rect 2789 12256 3036 12363
rect 2789 12219 2810 12256
rect 2789 12164 2809 12219
rect 2678 12104 2809 12164
rect 3030 12070 3036 12256
rect 3070 12070 3076 12546
rect 3030 12058 3076 12070
rect 3488 12546 3534 12558
rect 3488 12070 3494 12546
rect 3528 12359 3534 12546
rect 3583 12359 3661 14613
rect 3730 14422 3736 14613
rect 3770 14422 3776 14898
rect 3730 14410 3776 14422
rect 4188 14898 4234 14910
rect 4188 14422 4194 14898
rect 4228 14422 4234 14898
rect 4188 14410 4234 14422
rect 5810 14751 5852 14959
rect 5930 14943 7030 14949
rect 5930 14909 5942 14943
rect 7018 14909 7030 14943
rect 5930 14903 7030 14909
rect 5930 14801 7030 14807
rect 5930 14767 5942 14801
rect 7018 14767 7030 14801
rect 5930 14761 7030 14767
rect 7108 14753 7150 14959
rect 7376 14897 8476 14903
rect 7376 14863 7388 14897
rect 8464 14863 8476 14897
rect 7376 14857 8476 14863
rect 8714 14856 8749 14971
rect 8976 14954 8982 15082
rect 9016 14954 9022 15082
rect 8976 14942 9022 14954
rect 9304 15082 9350 15094
rect 9304 14954 9310 15082
rect 9344 14954 9350 15082
rect 9304 14942 9350 14954
rect 9667 15082 9713 15094
rect 9667 14954 9673 15082
rect 9707 14954 9713 15082
rect 9667 14942 9713 14954
rect 9995 15082 10041 15094
rect 9995 14954 10001 15082
rect 10035 14954 10041 15082
rect 10215 15079 10234 15162
rect 10269 15079 10287 15162
rect 10215 15063 10287 15079
rect 10385 15221 11737 15265
rect 10385 15129 10433 15221
rect 10511 15179 11611 15185
rect 10511 15145 10523 15179
rect 11599 15145 11611 15179
rect 10511 15139 11611 15145
rect 11689 15129 11737 15221
rect 10385 15117 10479 15129
rect 10385 15069 10439 15117
rect 10473 15069 10479 15117
rect 10385 15057 10479 15069
rect 11643 15117 11737 15129
rect 11643 15069 11649 15117
rect 11683 15069 11737 15117
rect 11643 15057 11737 15069
rect 11867 15459 11955 15471
rect 11867 15331 11915 15459
rect 11949 15331 11955 15459
rect 11867 15319 11955 15331
rect 13119 15459 13207 15471
rect 13119 15331 13125 15459
rect 13159 15331 13207 15459
rect 13119 15319 13207 15331
rect 11867 15111 11909 15319
rect 11987 15303 13087 15309
rect 11987 15269 11999 15303
rect 13075 15269 13087 15303
rect 11987 15263 13087 15269
rect 11987 15161 13087 15167
rect 11987 15127 11999 15161
rect 13075 15127 13087 15161
rect 11987 15121 13087 15127
rect 13165 15111 13207 15319
rect 18368 15242 18647 18292
rect 11867 15099 11955 15111
rect 10511 15041 11611 15047
rect 10511 15012 10523 15041
rect 9995 14942 10041 14954
rect 10268 15007 10523 15012
rect 11599 15007 11611 15041
rect 10268 15001 11611 15007
rect 10268 14971 10768 15001
rect 11867 14971 11915 15099
rect 11949 14971 11955 15099
rect 9063 14926 9263 14932
rect 9063 14892 9075 14926
rect 9251 14892 9263 14926
rect 9063 14886 9263 14892
rect 9754 14926 9954 14932
rect 9754 14892 9766 14926
rect 9942 14892 9954 14926
rect 9754 14886 9954 14892
rect 9126 14856 9196 14886
rect 7256 14835 7344 14847
rect 7256 14753 7304 14835
rect 7108 14751 7304 14753
rect 5810 14739 5898 14751
rect 5810 14611 5858 14739
rect 5892 14611 5898 14739
rect 5810 14599 5898 14611
rect 7062 14739 7304 14751
rect 7062 14611 7068 14739
rect 7102 14691 7304 14739
rect 7102 14643 7150 14691
rect 7256 14667 7304 14691
rect 7338 14667 7344 14835
rect 7256 14655 7344 14667
rect 8508 14835 8596 14847
rect 8508 14667 8514 14835
rect 8548 14667 8596 14835
rect 8714 14772 9196 14856
rect 9821 14856 9891 14886
rect 10268 14856 10303 14971
rect 11867 14959 11955 14971
rect 13119 15099 13207 15111
rect 13119 14971 13125 15099
rect 13159 14971 13207 15099
rect 13119 14959 13207 14971
rect 10541 14897 11641 14903
rect 10541 14863 10553 14897
rect 11629 14863 11641 14897
rect 10541 14857 11641 14863
rect 9126 14704 9196 14772
rect 9271 14829 9376 14851
rect 9271 14761 9291 14829
rect 9354 14761 9376 14829
rect 9271 14744 9376 14761
rect 9641 14829 9746 14851
rect 9641 14761 9663 14829
rect 9726 14761 9746 14829
rect 9641 14744 9746 14761
rect 9821 14772 10303 14856
rect 10421 14835 10509 14847
rect 9821 14704 9891 14772
rect 8508 14655 8596 14667
rect 9063 14698 9263 14704
rect 9063 14664 9075 14698
rect 9251 14664 9263 14698
rect 9063 14658 9263 14664
rect 9754 14698 9954 14704
rect 9754 14664 9766 14698
rect 9942 14664 9954 14698
rect 9754 14658 9954 14664
rect 10421 14667 10469 14835
rect 10503 14667 10509 14835
rect 7102 14611 7152 14643
rect 7062 14599 7152 14611
rect 5810 14391 5852 14599
rect 5930 14583 7030 14589
rect 5930 14549 5942 14583
rect 7018 14549 7030 14583
rect 5930 14543 7030 14549
rect 5930 14441 7030 14447
rect 5930 14407 5942 14441
rect 7018 14407 7030 14441
rect 5930 14401 7030 14407
rect 7108 14423 7152 14599
rect 7256 14561 7298 14655
rect 7376 14639 8476 14645
rect 7376 14605 7388 14639
rect 8464 14605 8476 14639
rect 7376 14599 8476 14605
rect 8554 14561 8596 14655
rect 10421 14655 10509 14667
rect 11673 14835 11761 14847
rect 11673 14667 11679 14835
rect 11713 14753 11761 14835
rect 11867 14753 11909 14959
rect 11987 14943 13087 14949
rect 11987 14909 11999 14943
rect 13075 14909 13087 14943
rect 11987 14903 13087 14909
rect 11987 14801 13087 14807
rect 11987 14767 11999 14801
rect 13075 14767 13087 14801
rect 11987 14761 13087 14767
rect 11713 14751 11909 14753
rect 13165 14751 13207 14959
rect 11713 14739 11955 14751
rect 11713 14691 11915 14739
rect 11713 14667 11761 14691
rect 11673 14655 11761 14667
rect 7256 14523 8596 14561
rect 7256 14423 7298 14523
rect 7376 14473 8476 14479
rect 7376 14439 7388 14473
rect 8464 14439 8476 14473
rect 7376 14433 8476 14439
rect 8554 14430 8596 14523
rect 8976 14636 9022 14648
rect 8976 14430 8982 14636
rect 8554 14423 8982 14430
rect 7108 14391 7150 14423
rect 5810 14379 5898 14391
rect 3786 14363 4178 14369
rect 3786 14329 3798 14363
rect 4166 14329 4178 14363
rect 3786 14207 4178 14329
rect 5810 14251 5858 14379
rect 5892 14251 5898 14379
rect 5810 14239 5898 14251
rect 7062 14379 7150 14391
rect 7062 14251 7068 14379
rect 7102 14369 7150 14379
rect 7256 14411 7344 14423
rect 7256 14369 7304 14411
rect 7102 14307 7304 14369
rect 7102 14251 7150 14307
rect 7062 14239 7150 14251
rect 7256 14243 7304 14307
rect 7338 14243 7344 14411
rect 7256 14231 7344 14243
rect 8508 14411 8982 14423
rect 8508 14243 8514 14411
rect 8548 14297 8982 14411
rect 8548 14243 8596 14297
rect 8976 14268 8982 14297
rect 9016 14268 9022 14636
rect 8976 14256 9022 14268
rect 9304 14636 9350 14648
rect 9304 14268 9310 14636
rect 9344 14268 9350 14636
rect 9304 14256 9350 14268
rect 9667 14636 9713 14648
rect 9667 14268 9673 14636
rect 9707 14268 9713 14636
rect 9667 14256 9713 14268
rect 9995 14636 10041 14648
rect 9995 14268 10001 14636
rect 10035 14430 10041 14636
rect 10421 14561 10463 14655
rect 10541 14639 11641 14645
rect 10541 14605 10553 14639
rect 11629 14605 11641 14639
rect 10541 14599 11641 14605
rect 11719 14561 11761 14655
rect 11867 14643 11915 14691
rect 10421 14523 11761 14561
rect 10421 14430 10463 14523
rect 10541 14473 11641 14479
rect 10541 14439 10553 14473
rect 11629 14439 11641 14473
rect 10541 14433 11641 14439
rect 10035 14423 10463 14430
rect 11719 14423 11761 14523
rect 11865 14611 11915 14643
rect 11949 14611 11955 14739
rect 11865 14599 11955 14611
rect 13119 14739 13207 14751
rect 13119 14611 13125 14739
rect 13159 14611 13207 14739
rect 13119 14599 13207 14611
rect 11865 14423 11909 14599
rect 11987 14583 13087 14589
rect 11987 14549 11999 14583
rect 13075 14549 13087 14583
rect 11987 14543 13087 14549
rect 10035 14411 10509 14423
rect 10035 14297 10469 14411
rect 10035 14268 10041 14297
rect 9995 14256 10041 14268
rect 8508 14231 8596 14243
rect 9063 14240 9263 14246
rect 3786 14173 3798 14207
rect 4166 14173 4178 14207
rect 5930 14223 7030 14229
rect 5930 14189 5942 14223
rect 7018 14189 7030 14223
rect 5930 14183 7030 14189
rect 7376 14215 8476 14221
rect 7376 14181 7388 14215
rect 8464 14181 8476 14215
rect 9063 14206 9075 14240
rect 9251 14206 9263 14240
rect 9063 14200 9263 14206
rect 9754 14240 9954 14246
rect 9754 14206 9766 14240
rect 9942 14206 9954 14240
rect 10421 14243 10469 14297
rect 10503 14243 10509 14411
rect 10421 14231 10509 14243
rect 11673 14411 11761 14423
rect 11673 14243 11679 14411
rect 11713 14369 11761 14411
rect 11867 14391 11909 14423
rect 11987 14441 13087 14447
rect 11987 14407 11999 14441
rect 13075 14407 13087 14441
rect 11987 14401 13087 14407
rect 13165 14391 13207 14599
rect 16133 14963 18647 15242
rect 16133 14550 16412 14963
rect 11867 14379 11955 14391
rect 11867 14369 11915 14379
rect 11713 14307 11915 14369
rect 11713 14243 11761 14307
rect 11673 14231 11761 14243
rect 11867 14251 11915 14307
rect 11949 14251 11955 14379
rect 11867 14239 11955 14251
rect 13119 14379 13207 14391
rect 13119 14251 13125 14379
rect 13159 14251 13207 14379
rect 13119 14239 13207 14251
rect 11987 14223 13087 14229
rect 9754 14200 9954 14206
rect 10541 14215 11641 14221
rect 7376 14175 8476 14181
rect 10541 14181 10553 14215
rect 11629 14181 11641 14215
rect 11987 14189 11999 14223
rect 13075 14189 13087 14223
rect 11987 14183 13087 14189
rect 10541 14175 11641 14181
rect 3786 14167 4178 14173
rect 3730 14114 3776 14126
rect 3730 13638 3736 14114
rect 3770 13638 3776 14114
rect 3730 13626 3776 13638
rect 4188 14114 4234 14126
rect 13596 14124 18558 14550
rect 4188 13638 4194 14114
rect 4228 13638 4234 14114
rect 8388 14058 8672 14059
rect 10345 14058 10629 14059
rect 8388 14041 9189 14058
rect 8388 13972 8416 14041
rect 8643 13972 9189 14041
rect 8388 13969 9189 13972
rect 8388 13959 8672 13969
rect 7125 13895 7330 13937
rect 6450 13861 8801 13895
rect 9130 13892 9189 13969
rect 9828 14041 10629 14058
rect 9828 13972 10374 14041
rect 10601 13972 10629 14041
rect 9828 13969 10629 13972
rect 9828 13892 9887 13969
rect 10345 13959 10629 13969
rect 11687 13895 11892 13937
rect 5930 13859 8801 13861
rect 5930 13855 7030 13859
rect 5930 13821 5942 13855
rect 7018 13821 7030 13855
rect 5930 13815 7030 13821
rect 7280 13855 8801 13859
rect 4188 13626 4234 13638
rect 5810 13793 5898 13805
rect 5810 13665 5858 13793
rect 5892 13665 5898 13793
rect 5810 13653 5898 13665
rect 7062 13793 7150 13805
rect 7062 13665 7068 13793
rect 7102 13665 7150 13793
rect 7062 13653 7150 13665
rect 3786 13579 4178 13585
rect 3786 13545 3798 13579
rect 4166 13545 4178 13579
rect 3786 13423 4178 13545
rect 3786 13389 3798 13423
rect 4166 13389 4178 13423
rect 3786 13383 4178 13389
rect 5810 13445 5852 13653
rect 5930 13637 7030 13643
rect 5930 13603 5942 13637
rect 7018 13603 7030 13637
rect 5930 13597 7030 13603
rect 5930 13495 7030 13501
rect 5930 13461 5942 13495
rect 7018 13461 7030 13495
rect 5930 13455 7030 13461
rect 7108 13445 7150 13653
rect 5810 13433 5898 13445
rect 3730 13330 3776 13342
rect 3730 12854 3736 13330
rect 3770 12854 3776 13330
rect 3730 12842 3776 12854
rect 4188 13330 4234 13342
rect 4188 12854 4194 13330
rect 4228 12854 4234 13330
rect 4188 12842 4234 12854
rect 5810 13305 5858 13433
rect 5892 13305 5898 13433
rect 5810 13293 5898 13305
rect 7062 13433 7150 13445
rect 7062 13305 7068 13433
rect 7102 13305 7150 13433
rect 7280 13761 7328 13855
rect 8733 13826 8801 13855
rect 9063 13886 9263 13892
rect 9063 13852 9075 13886
rect 9251 13852 9263 13886
rect 9063 13846 9263 13852
rect 9754 13886 9954 13892
rect 9754 13852 9766 13886
rect 9942 13852 9954 13886
rect 9754 13846 9954 13852
rect 10216 13861 12567 13895
rect 13597 13888 18558 14124
rect 13597 13886 18539 13888
rect 13599 13882 16256 13886
rect 10216 13859 13087 13861
rect 10216 13855 11737 13859
rect 8976 13826 9022 13836
rect 8733 13824 9022 13826
rect 7406 13811 8506 13817
rect 7406 13777 7418 13811
rect 8494 13777 8506 13811
rect 7406 13771 8506 13777
rect 8733 13766 8982 13824
rect 8733 13765 8801 13766
rect 7280 13749 7374 13761
rect 7280 13701 7334 13749
rect 7368 13701 7374 13749
rect 7280 13689 7374 13701
rect 8538 13749 8632 13761
rect 8538 13701 8544 13749
rect 8578 13701 8632 13749
rect 8538 13689 8632 13701
rect 7280 13599 7328 13689
rect 7406 13673 8506 13679
rect 7406 13639 7418 13673
rect 8494 13639 8506 13673
rect 7406 13633 8506 13639
rect 8584 13599 8632 13689
rect 8976 13696 8982 13766
rect 9016 13696 9022 13824
rect 8976 13684 9022 13696
rect 9304 13824 9350 13836
rect 9304 13696 9310 13824
rect 9344 13696 9350 13824
rect 9304 13684 9350 13696
rect 9667 13824 9713 13836
rect 9667 13696 9673 13824
rect 9707 13696 9713 13824
rect 9667 13684 9713 13696
rect 9995 13826 10041 13836
rect 10216 13826 10284 13855
rect 9995 13824 10284 13826
rect 9995 13696 10001 13824
rect 10035 13766 10284 13824
rect 10511 13811 11611 13817
rect 10511 13777 10523 13811
rect 11599 13777 11611 13811
rect 10511 13771 11611 13777
rect 10035 13696 10041 13766
rect 10216 13765 10284 13766
rect 11689 13761 11737 13855
rect 11987 13855 13087 13859
rect 11987 13821 11999 13855
rect 13075 13821 13087 13855
rect 11987 13815 13087 13821
rect 9995 13684 10041 13696
rect 10385 13749 10479 13761
rect 10385 13701 10439 13749
rect 10473 13701 10479 13749
rect 10385 13689 10479 13701
rect 11643 13749 11737 13761
rect 11643 13701 11649 13749
rect 11683 13701 11737 13749
rect 11643 13689 11737 13701
rect 9063 13668 9263 13674
rect 9063 13634 9075 13668
rect 9251 13634 9263 13668
rect 9063 13628 9263 13634
rect 9754 13668 9954 13674
rect 9754 13634 9766 13668
rect 9942 13634 9954 13668
rect 9754 13628 9954 13634
rect 7280 13555 8632 13599
rect 9143 13573 9187 13628
rect 7280 13463 7328 13555
rect 7406 13513 8506 13519
rect 7406 13479 7418 13513
rect 8494 13479 8506 13513
rect 7406 13473 8506 13479
rect 8584 13463 8632 13555
rect 7280 13451 7374 13463
rect 7280 13403 7334 13451
rect 7368 13403 7374 13451
rect 7280 13391 7374 13403
rect 8538 13451 8632 13463
rect 8538 13403 8544 13451
rect 8578 13403 8632 13451
rect 8538 13391 8632 13403
rect 8730 13528 9187 13573
rect 9249 13580 9436 13598
rect 9249 13528 9274 13580
rect 9372 13528 9436 13580
rect 8730 13496 8802 13528
rect 9249 13513 9436 13528
rect 9581 13580 9768 13598
rect 9581 13528 9645 13580
rect 9743 13528 9768 13580
rect 9830 13573 9874 13628
rect 10385 13599 10433 13689
rect 10511 13673 11611 13679
rect 10511 13639 10523 13673
rect 11599 13639 11611 13673
rect 10511 13633 11611 13639
rect 11689 13599 11737 13689
rect 9830 13528 10287 13573
rect 9581 13513 9768 13528
rect 8730 13413 8748 13496
rect 8783 13413 8802 13496
rect 10215 13496 10287 13528
rect 9063 13478 9263 13484
rect 9063 13444 9075 13478
rect 9251 13444 9263 13478
rect 9063 13438 9263 13444
rect 9754 13478 9954 13484
rect 9754 13444 9766 13478
rect 9942 13444 9954 13478
rect 9754 13438 9954 13444
rect 8730 13397 8802 13413
rect 8976 13416 9022 13428
rect 7406 13375 8506 13381
rect 7406 13341 7418 13375
rect 8494 13346 8506 13375
rect 8494 13341 8749 13346
rect 7406 13335 8749 13341
rect 8249 13305 8749 13335
rect 7062 13293 7150 13305
rect 5810 13085 5852 13293
rect 5930 13277 7030 13283
rect 5930 13243 5942 13277
rect 7018 13243 7030 13277
rect 5930 13237 7030 13243
rect 5930 13135 7030 13141
rect 5930 13101 5942 13135
rect 7018 13101 7030 13135
rect 5930 13095 7030 13101
rect 7108 13087 7150 13293
rect 7376 13231 8476 13237
rect 7376 13197 7388 13231
rect 8464 13197 8476 13231
rect 7376 13191 8476 13197
rect 8714 13190 8749 13305
rect 8976 13288 8982 13416
rect 9016 13288 9022 13416
rect 8976 13276 9022 13288
rect 9304 13416 9350 13428
rect 9304 13288 9310 13416
rect 9344 13288 9350 13416
rect 9304 13276 9350 13288
rect 9667 13416 9713 13428
rect 9667 13288 9673 13416
rect 9707 13288 9713 13416
rect 9667 13276 9713 13288
rect 9995 13416 10041 13428
rect 9995 13288 10001 13416
rect 10035 13288 10041 13416
rect 10215 13413 10234 13496
rect 10269 13413 10287 13496
rect 10215 13397 10287 13413
rect 10385 13555 11737 13599
rect 10385 13463 10433 13555
rect 10511 13513 11611 13519
rect 10511 13479 10523 13513
rect 11599 13479 11611 13513
rect 10511 13473 11611 13479
rect 11689 13463 11737 13555
rect 10385 13451 10479 13463
rect 10385 13403 10439 13451
rect 10473 13403 10479 13451
rect 10385 13391 10479 13403
rect 11643 13451 11737 13463
rect 11643 13403 11649 13451
rect 11683 13403 11737 13451
rect 11643 13391 11737 13403
rect 11867 13793 11955 13805
rect 11867 13665 11915 13793
rect 11949 13665 11955 13793
rect 11867 13653 11955 13665
rect 13119 13793 13207 13805
rect 13119 13665 13125 13793
rect 13159 13665 13207 13793
rect 13119 13653 13207 13665
rect 11867 13445 11909 13653
rect 11987 13637 13087 13643
rect 11987 13603 11999 13637
rect 13075 13603 13087 13637
rect 11987 13597 13087 13603
rect 11987 13495 13087 13501
rect 11987 13461 11999 13495
rect 13075 13461 13087 13495
rect 11987 13455 13087 13461
rect 13165 13445 13207 13653
rect 11867 13433 11955 13445
rect 10511 13375 11611 13381
rect 10511 13346 10523 13375
rect 9995 13276 10041 13288
rect 10268 13341 10523 13346
rect 11599 13341 11611 13375
rect 10268 13335 11611 13341
rect 10268 13305 10768 13335
rect 11867 13305 11915 13433
rect 11949 13305 11955 13433
rect 9063 13260 9263 13266
rect 9063 13226 9075 13260
rect 9251 13226 9263 13260
rect 9063 13220 9263 13226
rect 9754 13260 9954 13266
rect 9754 13226 9766 13260
rect 9942 13226 9954 13260
rect 9754 13220 9954 13226
rect 9126 13190 9196 13220
rect 7256 13169 7344 13181
rect 7256 13087 7304 13169
rect 7108 13085 7304 13087
rect 5810 13073 5898 13085
rect 5810 12945 5858 13073
rect 5892 12945 5898 13073
rect 5810 12933 5898 12945
rect 7062 13073 7304 13085
rect 7062 12945 7068 13073
rect 7102 13025 7304 13073
rect 7102 12977 7150 13025
rect 7256 13001 7304 13025
rect 7338 13001 7344 13169
rect 7256 12989 7344 13001
rect 8508 13169 8596 13181
rect 8508 13001 8514 13169
rect 8548 13001 8596 13169
rect 8714 13106 9196 13190
rect 9821 13190 9891 13220
rect 10268 13190 10303 13305
rect 11867 13293 11955 13305
rect 13119 13433 13207 13445
rect 13119 13305 13125 13433
rect 13159 13305 13207 13433
rect 13119 13293 13207 13305
rect 10541 13231 11641 13237
rect 10541 13197 10553 13231
rect 11629 13197 11641 13231
rect 10541 13191 11641 13197
rect 9126 13038 9196 13106
rect 9271 13163 9376 13185
rect 9271 13095 9291 13163
rect 9354 13095 9376 13163
rect 9271 13078 9376 13095
rect 9641 13163 9746 13185
rect 9641 13095 9663 13163
rect 9726 13095 9746 13163
rect 9641 13078 9746 13095
rect 9821 13106 10303 13190
rect 10421 13169 10509 13181
rect 9821 13038 9891 13106
rect 8508 12989 8596 13001
rect 9063 13032 9263 13038
rect 9063 12998 9075 13032
rect 9251 12998 9263 13032
rect 9063 12992 9263 12998
rect 9754 13032 9954 13038
rect 9754 12998 9766 13032
rect 9942 12998 9954 13032
rect 9754 12992 9954 12998
rect 10421 13001 10469 13169
rect 10503 13001 10509 13169
rect 7102 12945 7152 12977
rect 7062 12933 7152 12945
rect 3786 12795 4178 12801
rect 3786 12761 3798 12795
rect 4166 12761 4178 12795
rect 3786 12639 4178 12761
rect 3786 12605 3798 12639
rect 4166 12605 4178 12639
rect 3786 12599 4178 12605
rect 5810 12725 5852 12933
rect 5930 12917 7030 12923
rect 5930 12883 5942 12917
rect 7018 12883 7030 12917
rect 5930 12877 7030 12883
rect 5930 12775 7030 12781
rect 5930 12741 5942 12775
rect 7018 12741 7030 12775
rect 5930 12735 7030 12741
rect 7108 12757 7152 12933
rect 7256 12895 7298 12989
rect 7376 12973 8476 12979
rect 7376 12939 7388 12973
rect 8464 12939 8476 12973
rect 7376 12933 8476 12939
rect 8554 12895 8596 12989
rect 10421 12989 10509 13001
rect 11673 13169 11761 13181
rect 11673 13001 11679 13169
rect 11713 13087 11761 13169
rect 11867 13087 11909 13293
rect 11987 13277 13087 13283
rect 11987 13243 11999 13277
rect 13075 13243 13087 13277
rect 11987 13237 13087 13243
rect 11987 13135 13087 13141
rect 11987 13101 11999 13135
rect 13075 13101 13087 13135
rect 11987 13095 13087 13101
rect 11713 13085 11909 13087
rect 13165 13085 13207 13293
rect 11713 13073 11955 13085
rect 11713 13025 11915 13073
rect 11713 13001 11761 13025
rect 11673 12989 11761 13001
rect 7256 12857 8596 12895
rect 7256 12757 7298 12857
rect 7376 12807 8476 12813
rect 7376 12773 7388 12807
rect 8464 12773 8476 12807
rect 7376 12767 8476 12773
rect 8554 12764 8596 12857
rect 8976 12970 9022 12982
rect 8976 12764 8982 12970
rect 8554 12757 8982 12764
rect 7108 12725 7150 12757
rect 5810 12713 5898 12725
rect 5810 12585 5858 12713
rect 5892 12585 5898 12713
rect 5810 12573 5898 12585
rect 7062 12713 7150 12725
rect 7062 12585 7068 12713
rect 7102 12703 7150 12713
rect 7256 12745 7344 12757
rect 7256 12703 7304 12745
rect 7102 12641 7304 12703
rect 7102 12585 7150 12641
rect 7062 12573 7150 12585
rect 7256 12577 7304 12641
rect 7338 12577 7344 12745
rect 7256 12565 7344 12577
rect 8508 12745 8982 12757
rect 8508 12577 8514 12745
rect 8548 12631 8982 12745
rect 8548 12577 8596 12631
rect 8976 12602 8982 12631
rect 9016 12602 9022 12970
rect 8976 12590 9022 12602
rect 9304 12970 9350 12982
rect 9304 12602 9310 12970
rect 9344 12602 9350 12970
rect 9304 12590 9350 12602
rect 9667 12970 9713 12982
rect 9667 12602 9673 12970
rect 9707 12602 9713 12970
rect 9667 12590 9713 12602
rect 9995 12970 10041 12982
rect 9995 12602 10001 12970
rect 10035 12764 10041 12970
rect 10421 12895 10463 12989
rect 10541 12973 11641 12979
rect 10541 12939 10553 12973
rect 11629 12939 11641 12973
rect 10541 12933 11641 12939
rect 11719 12895 11761 12989
rect 11867 12977 11915 13025
rect 10421 12857 11761 12895
rect 10421 12764 10463 12857
rect 10541 12807 11641 12813
rect 10541 12773 10553 12807
rect 11629 12773 11641 12807
rect 10541 12767 11641 12773
rect 10035 12757 10463 12764
rect 11719 12757 11761 12857
rect 11865 12945 11915 12977
rect 11949 12945 11955 13073
rect 11865 12933 11955 12945
rect 13119 13073 13207 13085
rect 13119 12945 13125 13073
rect 13159 12945 13207 13073
rect 13119 12933 13207 12945
rect 11865 12757 11909 12933
rect 11987 12917 13087 12923
rect 11987 12883 11999 12917
rect 13075 12883 13087 12917
rect 11987 12877 13087 12883
rect 10035 12745 10509 12757
rect 10035 12631 10469 12745
rect 10035 12602 10041 12631
rect 9995 12590 10041 12602
rect 8508 12565 8596 12577
rect 9063 12574 9263 12580
rect 3730 12546 3776 12558
rect 3730 12359 3736 12546
rect 3528 12337 3736 12359
rect 3528 12273 3597 12337
rect 3653 12273 3736 12337
rect 3528 12252 3736 12273
rect 3528 12070 3534 12252
rect 3488 12058 3534 12070
rect 3730 12070 3736 12252
rect 3770 12070 3776 12546
rect 3730 12058 3776 12070
rect 4188 12546 4234 12558
rect 4188 12070 4194 12546
rect 4228 12070 4234 12546
rect 5930 12557 7030 12563
rect 5930 12523 5942 12557
rect 7018 12523 7030 12557
rect 5930 12517 7030 12523
rect 7376 12549 8476 12555
rect 7376 12515 7388 12549
rect 8464 12515 8476 12549
rect 9063 12540 9075 12574
rect 9251 12540 9263 12574
rect 9063 12534 9263 12540
rect 9754 12574 9954 12580
rect 9754 12540 9766 12574
rect 9942 12540 9954 12574
rect 10421 12577 10469 12631
rect 10503 12577 10509 12745
rect 10421 12565 10509 12577
rect 11673 12745 11761 12757
rect 11673 12577 11679 12745
rect 11713 12703 11761 12745
rect 11867 12725 11909 12757
rect 11987 12775 13087 12781
rect 11987 12741 11999 12775
rect 13075 12741 13087 12775
rect 11987 12735 13087 12741
rect 13165 12725 13207 12933
rect 11867 12713 11955 12725
rect 11867 12703 11915 12713
rect 11713 12641 11915 12703
rect 11713 12577 11761 12641
rect 11673 12565 11761 12577
rect 11867 12585 11915 12641
rect 11949 12585 11955 12713
rect 11867 12573 11955 12585
rect 13119 12713 13207 12725
rect 13119 12585 13125 12713
rect 13159 12585 13207 12713
rect 13119 12573 13207 12585
rect 11987 12557 13087 12563
rect 9754 12534 9954 12540
rect 10541 12549 11641 12555
rect 7376 12509 8476 12515
rect 10541 12515 10553 12549
rect 11629 12515 11641 12549
rect 11987 12523 11999 12557
rect 13075 12523 13087 12557
rect 11987 12517 13087 12523
rect 10541 12509 11641 12515
rect 8388 12392 8672 12393
rect 10345 12392 10629 12393
rect 8388 12375 9189 12392
rect 8388 12306 8416 12375
rect 8643 12306 9189 12375
rect 8388 12303 9189 12306
rect 8388 12293 8672 12303
rect 7125 12229 7330 12271
rect 6450 12195 8801 12229
rect 9130 12226 9189 12303
rect 9828 12375 10629 12392
rect 9828 12306 10374 12375
rect 10601 12306 10629 12375
rect 9828 12303 10629 12306
rect 9828 12226 9887 12303
rect 10345 12293 10629 12303
rect 11687 12229 11892 12271
rect 5930 12193 8801 12195
rect 5930 12189 7030 12193
rect 5930 12155 5942 12189
rect 7018 12155 7030 12189
rect 5930 12149 7030 12155
rect 7280 12189 8801 12193
rect 4188 12058 4234 12070
rect 5810 12127 5898 12139
rect 3086 12011 3478 12017
rect 783 11980 2169 11986
rect 783 11946 795 11980
rect 2157 11946 2169 11980
rect 783 11940 2169 11946
rect 3086 11977 3098 12011
rect 3466 11977 3478 12011
rect 727 11887 773 11899
rect 727 11877 733 11887
rect 499 11745 733 11877
rect 727 11735 733 11745
rect 767 11735 773 11887
rect 727 11723 773 11735
rect 2179 11887 2225 11899
rect 2179 11735 2185 11887
rect 2219 11735 2225 11887
rect 3086 11855 3478 11977
rect 3086 11821 3098 11855
rect 3466 11821 3478 11855
rect 3086 11815 3478 11821
rect 3786 12011 4178 12017
rect 3786 11977 3798 12011
rect 4166 11977 4178 12011
rect 3786 11855 4178 11977
rect 3786 11821 3798 11855
rect 4166 11821 4178 11855
rect 3786 11815 4178 11821
rect 5810 11999 5858 12127
rect 5892 11999 5898 12127
rect 5810 11987 5898 11999
rect 7062 12127 7150 12139
rect 7062 11999 7068 12127
rect 7102 11999 7150 12127
rect 7062 11987 7150 11999
rect 5810 11779 5852 11987
rect 5930 11971 7030 11977
rect 5930 11937 5942 11971
rect 7018 11937 7030 11971
rect 5930 11931 7030 11937
rect 5930 11829 7030 11835
rect 5930 11795 5942 11829
rect 7018 11795 7030 11829
rect 5930 11789 7030 11795
rect 7108 11779 7150 11987
rect 2179 11723 2225 11735
rect 2987 11762 3076 11774
rect 783 11676 2169 11682
rect 783 11642 795 11676
rect 2157 11642 2169 11676
rect 783 11636 2169 11642
rect 666 11510 925 11554
rect 666 11357 698 11510
rect 875 11357 925 11510
rect 666 11315 925 11357
rect 666 11084 819 11315
rect 2987 11286 3036 11762
rect 3070 11286 3076 11762
rect 2987 11274 3076 11286
rect 3488 11762 3534 11774
rect 3488 11286 3494 11762
rect 3528 11590 3534 11762
rect 3730 11762 3776 11774
rect 3730 11590 3736 11762
rect 3528 11582 3736 11590
rect 3528 11463 3598 11582
rect 3528 11286 3534 11463
rect 3488 11274 3534 11286
rect 3593 11300 3598 11463
rect 3653 11463 3736 11582
rect 3653 11300 3658 11463
rect 405 11078 951 11084
rect 405 11044 417 11078
rect 939 11044 951 11078
rect 405 11038 951 11044
rect 1399 11072 2247 11078
rect 1399 11038 1411 11072
rect 2179 11038 2247 11072
rect 1399 11032 2247 11038
rect 44 10985 395 10997
rect 44 10863 355 10985
rect 349 10323 355 10863
rect 389 10323 395 10985
rect 349 10311 395 10323
rect 961 10991 1007 10997
rect 2191 10991 2247 11032
rect 961 10985 1389 10991
rect 961 10323 967 10985
rect 1001 10979 1389 10985
rect 1001 10903 1349 10979
rect 1383 10903 1389 10979
rect 1001 10891 1389 10903
rect 2201 10979 2247 10991
rect 2987 10990 3030 11274
rect 3086 11227 3478 11233
rect 3086 11193 3098 11227
rect 3466 11193 3478 11227
rect 3086 11071 3478 11193
rect 3086 11037 3098 11071
rect 3466 11037 3478 11071
rect 3086 11031 3478 11037
rect 2201 10903 2207 10979
rect 2241 10903 2247 10979
rect 2201 10891 2247 10903
rect 1001 10323 1007 10891
rect 961 10311 1007 10323
rect 1134 10721 1171 10891
rect 2191 10850 2247 10891
rect 1399 10844 2247 10850
rect 1399 10810 1411 10844
rect 2179 10810 2247 10844
rect 1399 10804 2247 10810
rect 2934 10978 3076 10990
rect 2934 10907 3036 10978
rect 1134 10684 2193 10721
rect 405 10264 951 10270
rect 405 10230 417 10264
rect 939 10230 951 10264
rect 405 10224 951 10230
rect 1134 10049 1171 10684
rect 1325 10680 2193 10684
rect 1325 10646 1337 10680
rect 2181 10646 2193 10680
rect 1325 10640 2193 10646
rect 1269 10587 1315 10599
rect 1269 10137 1275 10587
rect 1309 10137 1315 10587
rect 1269 10125 1315 10137
rect 2203 10587 2249 10599
rect 2203 10137 2209 10587
rect 2243 10137 2249 10587
rect 2203 10125 2249 10137
rect 1325 10078 2193 10084
rect 1325 10049 1337 10078
rect 1134 10044 1337 10049
rect 2181 10044 2193 10078
rect 1134 10038 2193 10044
rect 1134 10007 2149 10038
rect 1060 9333 1551 9339
rect 1060 9299 1171 9333
rect 1539 9299 1551 9333
rect 1060 9293 1551 9299
rect 1859 9333 2251 9339
rect 1859 9299 1871 9333
rect 2239 9299 2251 9333
rect 1859 9293 2251 9299
rect 1060 9252 1159 9293
rect 1060 9240 1149 9252
rect 1060 8764 1109 9240
rect 1143 8764 1149 9240
rect 1060 8752 1149 8764
rect 1561 9240 1849 9252
rect 1561 8764 1567 9240
rect 1601 8764 1809 9240
rect 1843 8764 1849 9240
rect 1561 8752 1849 8764
rect 2261 9240 2307 9252
rect 2261 8764 2267 9240
rect 2301 8764 2307 9240
rect 2261 8752 2307 8764
rect 2376 9116 2814 9166
rect 1060 8711 1159 8752
rect 1060 8705 1551 8711
rect 1060 8671 1171 8705
rect 1539 8671 1551 8705
rect 1060 8549 1551 8671
rect 1060 8515 1171 8549
rect 1539 8515 1551 8549
rect 1060 8509 1551 8515
rect 1660 8665 1803 8752
rect 1859 8705 2251 8711
rect 1859 8671 1871 8705
rect 2239 8671 2251 8705
rect 1859 8665 2251 8671
rect 1660 8555 2251 8665
rect 1060 8468 1159 8509
rect 1660 8468 1803 8555
rect 1859 8549 2251 8555
rect 1859 8515 1871 8549
rect 2239 8515 2251 8549
rect 1859 8509 2251 8515
rect 2376 8504 2420 9116
rect 2762 8504 2814 9116
rect 2934 8995 2954 10907
rect 3006 10502 3036 10907
rect 3070 10502 3076 10978
rect 3006 10490 3076 10502
rect 3488 10978 3534 10990
rect 3488 10502 3494 10978
rect 3528 10806 3534 10978
rect 3593 10806 3658 11300
rect 3730 11286 3736 11463
rect 3770 11286 3776 11762
rect 3730 11274 3776 11286
rect 4188 11762 4234 11774
rect 4188 11286 4194 11762
rect 4228 11286 4234 11762
rect 4188 11274 4234 11286
rect 5810 11767 5898 11779
rect 5810 11639 5858 11767
rect 5892 11639 5898 11767
rect 5810 11627 5898 11639
rect 7062 11767 7150 11779
rect 7062 11639 7068 11767
rect 7102 11639 7150 11767
rect 7280 12095 7328 12189
rect 8733 12160 8801 12189
rect 9063 12220 9263 12226
rect 9063 12186 9075 12220
rect 9251 12186 9263 12220
rect 9063 12180 9263 12186
rect 9754 12220 9954 12226
rect 9754 12186 9766 12220
rect 9942 12186 9954 12220
rect 9754 12180 9954 12186
rect 10216 12195 12567 12229
rect 10216 12193 13087 12195
rect 10216 12189 11737 12193
rect 8976 12160 9022 12170
rect 8733 12158 9022 12160
rect 7406 12145 8506 12151
rect 7406 12111 7418 12145
rect 8494 12111 8506 12145
rect 7406 12105 8506 12111
rect 8733 12100 8982 12158
rect 8733 12099 8801 12100
rect 7280 12083 7374 12095
rect 7280 12035 7334 12083
rect 7368 12035 7374 12083
rect 7280 12023 7374 12035
rect 8538 12083 8632 12095
rect 8538 12035 8544 12083
rect 8578 12035 8632 12083
rect 8538 12023 8632 12035
rect 7280 11933 7328 12023
rect 7406 12007 8506 12013
rect 7406 11973 7418 12007
rect 8494 11973 8506 12007
rect 7406 11967 8506 11973
rect 8584 11933 8632 12023
rect 8976 12030 8982 12100
rect 9016 12030 9022 12158
rect 8976 12018 9022 12030
rect 9304 12158 9350 12170
rect 9304 12030 9310 12158
rect 9344 12030 9350 12158
rect 9304 12018 9350 12030
rect 9667 12158 9713 12170
rect 9667 12030 9673 12158
rect 9707 12030 9713 12158
rect 9667 12018 9713 12030
rect 9995 12160 10041 12170
rect 10216 12160 10284 12189
rect 9995 12158 10284 12160
rect 9995 12030 10001 12158
rect 10035 12100 10284 12158
rect 10511 12145 11611 12151
rect 10511 12111 10523 12145
rect 11599 12111 11611 12145
rect 10511 12105 11611 12111
rect 10035 12030 10041 12100
rect 10216 12099 10284 12100
rect 11689 12095 11737 12189
rect 11987 12189 13087 12193
rect 11987 12155 11999 12189
rect 13075 12155 13087 12189
rect 11987 12149 13087 12155
rect 9995 12018 10041 12030
rect 10385 12083 10479 12095
rect 10385 12035 10439 12083
rect 10473 12035 10479 12083
rect 10385 12023 10479 12035
rect 11643 12083 11737 12095
rect 11643 12035 11649 12083
rect 11683 12035 11737 12083
rect 11643 12023 11737 12035
rect 9063 12002 9263 12008
rect 9063 11968 9075 12002
rect 9251 11968 9263 12002
rect 9063 11962 9263 11968
rect 9754 12002 9954 12008
rect 9754 11968 9766 12002
rect 9942 11968 9954 12002
rect 9754 11962 9954 11968
rect 7280 11889 8632 11933
rect 9143 11907 9187 11962
rect 7280 11797 7328 11889
rect 7406 11847 8506 11853
rect 7406 11813 7418 11847
rect 8494 11813 8506 11847
rect 7406 11807 8506 11813
rect 8584 11797 8632 11889
rect 7280 11785 7374 11797
rect 7280 11737 7334 11785
rect 7368 11737 7374 11785
rect 7280 11725 7374 11737
rect 8538 11785 8632 11797
rect 8538 11737 8544 11785
rect 8578 11737 8632 11785
rect 8538 11725 8632 11737
rect 8730 11862 9187 11907
rect 9249 11914 9436 11932
rect 9249 11862 9274 11914
rect 9372 11862 9436 11914
rect 8730 11830 8802 11862
rect 9249 11847 9436 11862
rect 9581 11914 9768 11932
rect 9581 11862 9645 11914
rect 9743 11862 9768 11914
rect 9830 11907 9874 11962
rect 10385 11933 10433 12023
rect 10511 12007 11611 12013
rect 10511 11973 10523 12007
rect 11599 11973 11611 12007
rect 10511 11967 11611 11973
rect 11689 11933 11737 12023
rect 9830 11862 10287 11907
rect 9581 11847 9768 11862
rect 8730 11747 8748 11830
rect 8783 11747 8802 11830
rect 10215 11830 10287 11862
rect 9063 11812 9263 11818
rect 9063 11778 9075 11812
rect 9251 11778 9263 11812
rect 9063 11772 9263 11778
rect 9754 11812 9954 11818
rect 9754 11778 9766 11812
rect 9942 11778 9954 11812
rect 9754 11772 9954 11778
rect 8730 11731 8802 11747
rect 8976 11750 9022 11762
rect 7406 11709 8506 11715
rect 7406 11675 7418 11709
rect 8494 11680 8506 11709
rect 8494 11675 8749 11680
rect 7406 11669 8749 11675
rect 8249 11639 8749 11669
rect 7062 11627 7150 11639
rect 5810 11419 5852 11627
rect 5930 11611 7030 11617
rect 5930 11577 5942 11611
rect 7018 11577 7030 11611
rect 5930 11571 7030 11577
rect 5930 11469 7030 11475
rect 5930 11435 5942 11469
rect 7018 11435 7030 11469
rect 5930 11429 7030 11435
rect 7108 11421 7150 11627
rect 7376 11565 8476 11571
rect 7376 11531 7388 11565
rect 8464 11531 8476 11565
rect 7376 11525 8476 11531
rect 8714 11524 8749 11639
rect 8976 11622 8982 11750
rect 9016 11622 9022 11750
rect 8976 11610 9022 11622
rect 9304 11750 9350 11762
rect 9304 11622 9310 11750
rect 9344 11622 9350 11750
rect 9304 11610 9350 11622
rect 9667 11750 9713 11762
rect 9667 11622 9673 11750
rect 9707 11622 9713 11750
rect 9667 11610 9713 11622
rect 9995 11750 10041 11762
rect 9995 11622 10001 11750
rect 10035 11622 10041 11750
rect 10215 11747 10234 11830
rect 10269 11747 10287 11830
rect 10215 11731 10287 11747
rect 10385 11889 11737 11933
rect 10385 11797 10433 11889
rect 10511 11847 11611 11853
rect 10511 11813 10523 11847
rect 11599 11813 11611 11847
rect 10511 11807 11611 11813
rect 11689 11797 11737 11889
rect 10385 11785 10479 11797
rect 10385 11737 10439 11785
rect 10473 11737 10479 11785
rect 10385 11725 10479 11737
rect 11643 11785 11737 11797
rect 11643 11737 11649 11785
rect 11683 11737 11737 11785
rect 11643 11725 11737 11737
rect 11867 12127 11955 12139
rect 11867 11999 11915 12127
rect 11949 11999 11955 12127
rect 11867 11987 11955 11999
rect 13119 12127 13207 12139
rect 13119 11999 13125 12127
rect 13159 11999 13207 12127
rect 13119 11987 13207 11999
rect 11867 11779 11909 11987
rect 11987 11971 13087 11977
rect 11987 11937 11999 11971
rect 13075 11937 13087 11971
rect 11987 11931 13087 11937
rect 11987 11829 13087 11835
rect 11987 11795 11999 11829
rect 13075 11795 13087 11829
rect 11987 11789 13087 11795
rect 13165 11779 13207 11987
rect 11867 11767 11955 11779
rect 10511 11709 11611 11715
rect 10511 11680 10523 11709
rect 9995 11610 10041 11622
rect 10268 11675 10523 11680
rect 11599 11675 11611 11709
rect 10268 11669 11611 11675
rect 10268 11639 10768 11669
rect 11867 11639 11915 11767
rect 11949 11639 11955 11767
rect 9063 11594 9263 11600
rect 9063 11560 9075 11594
rect 9251 11560 9263 11594
rect 9063 11554 9263 11560
rect 9754 11594 9954 11600
rect 9754 11560 9766 11594
rect 9942 11560 9954 11594
rect 9754 11554 9954 11560
rect 9126 11524 9196 11554
rect 7256 11503 7344 11515
rect 7256 11421 7304 11503
rect 7108 11419 7304 11421
rect 5810 11407 5898 11419
rect 5810 11279 5858 11407
rect 5892 11279 5898 11407
rect 5810 11267 5898 11279
rect 7062 11407 7304 11419
rect 7062 11279 7068 11407
rect 7102 11359 7304 11407
rect 7102 11311 7150 11359
rect 7256 11335 7304 11359
rect 7338 11335 7344 11503
rect 7256 11323 7344 11335
rect 8508 11503 8596 11515
rect 8508 11335 8514 11503
rect 8548 11335 8596 11503
rect 8714 11440 9196 11524
rect 9821 11524 9891 11554
rect 10268 11524 10303 11639
rect 11867 11627 11955 11639
rect 13119 11767 13207 11779
rect 13119 11639 13125 11767
rect 13159 11639 13207 11767
rect 13119 11627 13207 11639
rect 10541 11565 11641 11571
rect 10541 11531 10553 11565
rect 11629 11531 11641 11565
rect 10541 11525 11641 11531
rect 9126 11372 9196 11440
rect 9271 11497 9376 11519
rect 9271 11429 9291 11497
rect 9354 11429 9376 11497
rect 9271 11412 9376 11429
rect 9641 11497 9746 11519
rect 9641 11429 9663 11497
rect 9726 11429 9746 11497
rect 9641 11412 9746 11429
rect 9821 11440 10303 11524
rect 10421 11503 10509 11515
rect 9821 11372 9891 11440
rect 8508 11323 8596 11335
rect 9063 11366 9263 11372
rect 9063 11332 9075 11366
rect 9251 11332 9263 11366
rect 9063 11326 9263 11332
rect 9754 11366 9954 11372
rect 9754 11332 9766 11366
rect 9942 11332 9954 11366
rect 9754 11326 9954 11332
rect 10421 11335 10469 11503
rect 10503 11335 10509 11503
rect 7102 11279 7152 11311
rect 7062 11267 7152 11279
rect 3786 11227 4178 11233
rect 3786 11193 3798 11227
rect 4166 11193 4178 11227
rect 3786 11071 4178 11193
rect 3786 11037 3798 11071
rect 4166 11037 4178 11071
rect 3786 11031 4178 11037
rect 5810 11059 5852 11267
rect 5930 11251 7030 11257
rect 5930 11217 5942 11251
rect 7018 11217 7030 11251
rect 5930 11211 7030 11217
rect 5930 11109 7030 11115
rect 5930 11075 5942 11109
rect 7018 11075 7030 11109
rect 5930 11069 7030 11075
rect 7108 11091 7152 11267
rect 7256 11229 7298 11323
rect 7376 11307 8476 11313
rect 7376 11273 7388 11307
rect 8464 11273 8476 11307
rect 7376 11267 8476 11273
rect 8554 11229 8596 11323
rect 10421 11323 10509 11335
rect 11673 11503 11761 11515
rect 11673 11335 11679 11503
rect 11713 11421 11761 11503
rect 11867 11421 11909 11627
rect 11987 11611 13087 11617
rect 11987 11577 11999 11611
rect 13075 11577 13087 11611
rect 11987 11571 13087 11577
rect 11987 11469 13087 11475
rect 11987 11435 11999 11469
rect 13075 11435 13087 11469
rect 11987 11429 13087 11435
rect 11713 11419 11909 11421
rect 13165 11419 13207 11627
rect 11713 11407 11955 11419
rect 11713 11359 11915 11407
rect 11713 11335 11761 11359
rect 11673 11323 11761 11335
rect 7256 11191 8596 11229
rect 7256 11091 7298 11191
rect 7376 11141 8476 11147
rect 7376 11107 7388 11141
rect 8464 11107 8476 11141
rect 7376 11101 8476 11107
rect 8554 11098 8596 11191
rect 8976 11304 9022 11316
rect 8976 11098 8982 11304
rect 8554 11091 8982 11098
rect 7108 11059 7150 11091
rect 5810 11047 5898 11059
rect 3730 10978 3776 10990
rect 3730 10806 3736 10978
rect 3528 10679 3736 10806
rect 3528 10502 3534 10679
rect 3488 10490 3534 10502
rect 3006 10206 3030 10490
rect 3086 10443 3478 10449
rect 3086 10409 3098 10443
rect 3466 10409 3478 10443
rect 3086 10287 3478 10409
rect 3086 10253 3098 10287
rect 3466 10253 3478 10287
rect 3086 10247 3478 10253
rect 3006 10194 3076 10206
rect 3006 9718 3036 10194
rect 3070 9718 3076 10194
rect 3006 9706 3076 9718
rect 3488 10194 3534 10206
rect 3488 9718 3494 10194
rect 3528 10022 3534 10194
rect 3593 10022 3658 10679
rect 3730 10502 3736 10679
rect 3770 10502 3776 10978
rect 3730 10490 3776 10502
rect 4188 10978 4234 10990
rect 4188 10502 4194 10978
rect 4228 10502 4234 10978
rect 5810 10919 5858 11047
rect 5892 10919 5898 11047
rect 5810 10907 5898 10919
rect 7062 11047 7150 11059
rect 7062 10919 7068 11047
rect 7102 11037 7150 11047
rect 7256 11079 7344 11091
rect 7256 11037 7304 11079
rect 7102 10975 7304 11037
rect 7102 10919 7150 10975
rect 7062 10907 7150 10919
rect 7256 10911 7304 10975
rect 7338 10911 7344 11079
rect 7256 10899 7344 10911
rect 8508 11079 8982 11091
rect 8508 10911 8514 11079
rect 8548 10965 8982 11079
rect 8548 10911 8596 10965
rect 8976 10936 8982 10965
rect 9016 10936 9022 11304
rect 8976 10924 9022 10936
rect 9304 11304 9350 11316
rect 9304 10936 9310 11304
rect 9344 10936 9350 11304
rect 9304 10924 9350 10936
rect 9667 11304 9713 11316
rect 9667 10936 9673 11304
rect 9707 10936 9713 11304
rect 9667 10924 9713 10936
rect 9995 11304 10041 11316
rect 9995 10936 10001 11304
rect 10035 11098 10041 11304
rect 10421 11229 10463 11323
rect 10541 11307 11641 11313
rect 10541 11273 10553 11307
rect 11629 11273 11641 11307
rect 10541 11267 11641 11273
rect 11719 11229 11761 11323
rect 11867 11311 11915 11359
rect 10421 11191 11761 11229
rect 10421 11098 10463 11191
rect 10541 11141 11641 11147
rect 10541 11107 10553 11141
rect 11629 11107 11641 11141
rect 10541 11101 11641 11107
rect 10035 11091 10463 11098
rect 11719 11091 11761 11191
rect 11865 11279 11915 11311
rect 11949 11279 11955 11407
rect 11865 11267 11955 11279
rect 13119 11407 13207 11419
rect 13119 11279 13125 11407
rect 13159 11279 13207 11407
rect 13119 11267 13207 11279
rect 11865 11091 11909 11267
rect 11987 11251 13087 11257
rect 11987 11217 11999 11251
rect 13075 11217 13087 11251
rect 11987 11211 13087 11217
rect 10035 11079 10509 11091
rect 10035 10965 10469 11079
rect 10035 10936 10041 10965
rect 9995 10924 10041 10936
rect 8508 10899 8596 10911
rect 9063 10908 9263 10914
rect 5930 10891 7030 10897
rect 5930 10857 5942 10891
rect 7018 10857 7030 10891
rect 5930 10851 7030 10857
rect 7376 10883 8476 10889
rect 7376 10849 7388 10883
rect 8464 10849 8476 10883
rect 9063 10874 9075 10908
rect 9251 10874 9263 10908
rect 9063 10868 9263 10874
rect 9754 10908 9954 10914
rect 9754 10874 9766 10908
rect 9942 10874 9954 10908
rect 10421 10911 10469 10965
rect 10503 10911 10509 11079
rect 10421 10899 10509 10911
rect 11673 11079 11761 11091
rect 11673 10911 11679 11079
rect 11713 11037 11761 11079
rect 11867 11059 11909 11091
rect 11987 11109 13087 11115
rect 11987 11075 11999 11109
rect 13075 11075 13087 11109
rect 11987 11069 13087 11075
rect 13165 11059 13207 11267
rect 11867 11047 11955 11059
rect 11867 11037 11915 11047
rect 11713 10975 11915 11037
rect 11713 10911 11761 10975
rect 11673 10899 11761 10911
rect 11867 10919 11915 10975
rect 11949 10919 11955 11047
rect 11867 10907 11955 10919
rect 13119 11047 13207 11059
rect 13119 10919 13125 11047
rect 13159 10919 13207 11047
rect 13119 10907 13207 10919
rect 11987 10891 13087 10897
rect 9754 10868 9954 10874
rect 10541 10883 11641 10889
rect 7376 10843 8476 10849
rect 10541 10849 10553 10883
rect 11629 10849 11641 10883
rect 11987 10857 11999 10891
rect 13075 10857 13087 10891
rect 11987 10851 13087 10857
rect 10541 10843 11641 10849
rect 8388 10726 8672 10727
rect 10345 10726 10629 10727
rect 8388 10709 9189 10726
rect 8388 10640 8416 10709
rect 8643 10640 9189 10709
rect 8388 10637 9189 10640
rect 8388 10627 8672 10637
rect 7125 10563 7330 10605
rect 6450 10529 8801 10563
rect 9130 10560 9189 10637
rect 9828 10709 10629 10726
rect 9828 10640 10374 10709
rect 10601 10640 10629 10709
rect 9828 10637 10629 10640
rect 9828 10560 9887 10637
rect 10345 10627 10629 10637
rect 11687 10563 11892 10605
rect 4188 10490 4234 10502
rect 5930 10527 8801 10529
rect 5930 10523 7030 10527
rect 5930 10489 5942 10523
rect 7018 10489 7030 10523
rect 5930 10483 7030 10489
rect 7280 10523 8801 10527
rect 5810 10461 5898 10473
rect 3786 10443 4178 10449
rect 3786 10409 3798 10443
rect 4166 10409 4178 10443
rect 3786 10287 4178 10409
rect 3786 10253 3798 10287
rect 4166 10253 4178 10287
rect 3786 10247 4178 10253
rect 5810 10333 5858 10461
rect 5892 10333 5898 10461
rect 5810 10321 5898 10333
rect 7062 10461 7150 10473
rect 7062 10333 7068 10461
rect 7102 10333 7150 10461
rect 7062 10321 7150 10333
rect 3730 10194 3776 10206
rect 3730 10022 3736 10194
rect 3528 9895 3736 10022
rect 3528 9718 3534 9895
rect 3488 9706 3534 9718
rect 3006 9422 3030 9706
rect 3086 9659 3478 9665
rect 3086 9625 3098 9659
rect 3466 9625 3478 9659
rect 3086 9503 3478 9625
rect 3086 9469 3098 9503
rect 3466 9469 3478 9503
rect 3086 9463 3478 9469
rect 3006 9410 3076 9422
rect 3006 8995 3036 9410
rect 2934 8934 3036 8995
rect 3070 8934 3076 9410
rect 2934 8922 3076 8934
rect 3488 9410 3534 9422
rect 3488 8934 3494 9410
rect 3528 9238 3534 9410
rect 3593 9238 3658 9895
rect 3730 9718 3736 9895
rect 3770 9718 3776 10194
rect 3730 9706 3776 9718
rect 4188 10194 4234 10206
rect 4188 9718 4194 10194
rect 4228 9718 4234 10194
rect 5810 10113 5852 10321
rect 5930 10305 7030 10311
rect 5930 10271 5942 10305
rect 7018 10271 7030 10305
rect 5930 10265 7030 10271
rect 5930 10163 7030 10169
rect 5930 10129 5942 10163
rect 7018 10129 7030 10163
rect 5930 10123 7030 10129
rect 7108 10113 7150 10321
rect 5810 10101 5898 10113
rect 5810 9973 5858 10101
rect 5892 9973 5898 10101
rect 5810 9961 5898 9973
rect 7062 10101 7150 10113
rect 7062 9973 7068 10101
rect 7102 9973 7150 10101
rect 7280 10429 7328 10523
rect 8733 10494 8801 10523
rect 9063 10554 9263 10560
rect 9063 10520 9075 10554
rect 9251 10520 9263 10554
rect 9063 10514 9263 10520
rect 9754 10554 9954 10560
rect 9754 10520 9766 10554
rect 9942 10520 9954 10554
rect 9754 10514 9954 10520
rect 10216 10529 12567 10563
rect 10216 10527 13087 10529
rect 10216 10523 11737 10527
rect 8976 10494 9022 10504
rect 8733 10492 9022 10494
rect 7406 10479 8506 10485
rect 7406 10445 7418 10479
rect 8494 10445 8506 10479
rect 7406 10439 8506 10445
rect 8733 10434 8982 10492
rect 8733 10433 8801 10434
rect 7280 10417 7374 10429
rect 7280 10369 7334 10417
rect 7368 10369 7374 10417
rect 7280 10357 7374 10369
rect 8538 10417 8632 10429
rect 8538 10369 8544 10417
rect 8578 10369 8632 10417
rect 8538 10357 8632 10369
rect 7280 10267 7328 10357
rect 7406 10341 8506 10347
rect 7406 10307 7418 10341
rect 8494 10307 8506 10341
rect 7406 10301 8506 10307
rect 8584 10267 8632 10357
rect 8976 10364 8982 10434
rect 9016 10364 9022 10492
rect 8976 10352 9022 10364
rect 9304 10492 9350 10504
rect 9304 10364 9310 10492
rect 9344 10364 9350 10492
rect 9304 10352 9350 10364
rect 9667 10492 9713 10504
rect 9667 10364 9673 10492
rect 9707 10364 9713 10492
rect 9667 10352 9713 10364
rect 9995 10494 10041 10504
rect 10216 10494 10284 10523
rect 9995 10492 10284 10494
rect 9995 10364 10001 10492
rect 10035 10434 10284 10492
rect 10511 10479 11611 10485
rect 10511 10445 10523 10479
rect 11599 10445 11611 10479
rect 10511 10439 11611 10445
rect 10035 10364 10041 10434
rect 10216 10433 10284 10434
rect 11689 10429 11737 10523
rect 11987 10523 13087 10527
rect 11987 10489 11999 10523
rect 13075 10489 13087 10523
rect 11987 10483 13087 10489
rect 9995 10352 10041 10364
rect 10385 10417 10479 10429
rect 10385 10369 10439 10417
rect 10473 10369 10479 10417
rect 10385 10357 10479 10369
rect 11643 10417 11737 10429
rect 11643 10369 11649 10417
rect 11683 10369 11737 10417
rect 11643 10357 11737 10369
rect 9063 10336 9263 10342
rect 9063 10302 9075 10336
rect 9251 10302 9263 10336
rect 9063 10296 9263 10302
rect 9754 10336 9954 10342
rect 9754 10302 9766 10336
rect 9942 10302 9954 10336
rect 9754 10296 9954 10302
rect 7280 10223 8632 10267
rect 9143 10241 9187 10296
rect 7280 10131 7328 10223
rect 7406 10181 8506 10187
rect 7406 10147 7418 10181
rect 8494 10147 8506 10181
rect 7406 10141 8506 10147
rect 8584 10131 8632 10223
rect 7280 10119 7374 10131
rect 7280 10071 7334 10119
rect 7368 10071 7374 10119
rect 7280 10059 7374 10071
rect 8538 10119 8632 10131
rect 8538 10071 8544 10119
rect 8578 10071 8632 10119
rect 8538 10059 8632 10071
rect 8730 10196 9187 10241
rect 9249 10248 9436 10266
rect 9249 10196 9274 10248
rect 9372 10196 9436 10248
rect 8730 10164 8802 10196
rect 9249 10181 9436 10196
rect 9581 10248 9768 10266
rect 9581 10196 9645 10248
rect 9743 10196 9768 10248
rect 9830 10241 9874 10296
rect 10385 10267 10433 10357
rect 10511 10341 11611 10347
rect 10511 10307 10523 10341
rect 11599 10307 11611 10341
rect 10511 10301 11611 10307
rect 11689 10267 11737 10357
rect 9830 10196 10287 10241
rect 9581 10181 9768 10196
rect 8730 10081 8748 10164
rect 8783 10081 8802 10164
rect 10215 10164 10287 10196
rect 9063 10146 9263 10152
rect 9063 10112 9075 10146
rect 9251 10112 9263 10146
rect 9063 10106 9263 10112
rect 9754 10146 9954 10152
rect 9754 10112 9766 10146
rect 9942 10112 9954 10146
rect 9754 10106 9954 10112
rect 8730 10065 8802 10081
rect 8976 10084 9022 10096
rect 7406 10043 8506 10049
rect 7406 10009 7418 10043
rect 8494 10014 8506 10043
rect 8494 10009 8749 10014
rect 7406 10003 8749 10009
rect 8249 9973 8749 10003
rect 7062 9961 7150 9973
rect 4188 9706 4234 9718
rect 4766 9676 5354 9772
rect 3786 9659 4178 9665
rect 3786 9625 3798 9659
rect 4166 9625 4178 9659
rect 3786 9503 4178 9625
rect 3786 9469 3798 9503
rect 4166 9469 4178 9503
rect 3786 9463 4178 9469
rect 3730 9410 3776 9422
rect 3730 9238 3736 9410
rect 3528 9111 3736 9238
rect 3528 8934 3534 9111
rect 3488 8922 3534 8934
rect 1060 8456 1149 8468
rect 1060 7980 1109 8456
rect 1143 7980 1149 8456
rect 1060 7968 1149 7980
rect 1561 8456 1849 8468
rect 1561 7980 1567 8456
rect 1601 7980 1809 8456
rect 1843 7980 1849 8456
rect 1561 7968 1849 7980
rect 2261 8456 2307 8468
rect 2261 7980 2267 8456
rect 2301 7980 2307 8456
rect 2376 8454 2814 8504
rect 2987 8638 3030 8922
rect 3086 8875 3478 8881
rect 3086 8841 3098 8875
rect 3466 8841 3478 8875
rect 3086 8719 3478 8841
rect 3086 8685 3098 8719
rect 3466 8685 3478 8719
rect 3086 8679 3478 8685
rect 2987 8626 3076 8638
rect 2987 8150 3036 8626
rect 3070 8150 3076 8626
rect 2987 8138 3076 8150
rect 3488 8626 3534 8638
rect 3488 8150 3494 8626
rect 3528 8454 3534 8626
rect 3593 8454 3658 9111
rect 3730 8934 3736 9111
rect 3770 8934 3776 9410
rect 3730 8922 3776 8934
rect 4188 9410 4234 9422
rect 4188 8934 4194 9410
rect 4228 8934 4234 9410
rect 4188 8922 4234 8934
rect 3786 8875 4178 8881
rect 3786 8841 3798 8875
rect 4166 8841 4178 8875
rect 3786 8827 4178 8841
rect 3786 8735 3874 8827
rect 4110 8735 4178 8827
rect 3786 8719 4178 8735
rect 3786 8685 3798 8719
rect 4166 8685 4178 8719
rect 3786 8679 4178 8685
rect 3730 8626 3776 8638
rect 3730 8454 3736 8626
rect 3528 8327 3736 8454
rect 3528 8150 3534 8327
rect 3488 8138 3534 8150
rect 3730 8150 3736 8327
rect 3770 8150 3776 8626
rect 3730 8138 3776 8150
rect 4188 8626 4234 8638
rect 4188 8150 4194 8626
rect 4228 8150 4234 8626
rect 4188 8138 4234 8150
rect 3086 8091 3478 8097
rect 3086 8057 3098 8091
rect 3466 8057 3478 8091
rect 3086 8052 3478 8057
rect 2261 7968 2307 7980
rect 2696 8051 3478 8052
rect 3786 8091 4178 8097
rect 3786 8057 3798 8091
rect 4166 8057 4178 8091
rect 3786 8051 4178 8057
rect 2696 8008 3477 8051
rect 1060 7927 1159 7968
rect 1060 7921 1551 7927
rect -347 7832 116 7893
rect 1060 7887 1171 7921
rect 1539 7887 1551 7921
rect 1060 7881 1551 7887
rect 1859 7921 2251 7927
rect 1859 7887 1871 7921
rect 2239 7887 2251 7921
rect 1859 7881 2251 7887
rect -347 7595 -291 7832
rect 59 7759 116 7832
rect 1066 7759 1167 7881
rect 59 7695 1167 7759
rect 2696 7695 2765 8008
rect 3086 7935 3478 7941
rect 3086 7901 3098 7935
rect 3466 7901 3478 7935
rect 3086 7895 3478 7901
rect 3786 7935 4178 7941
rect 3786 7901 3798 7935
rect 4166 7901 4178 7935
rect 3786 7895 4178 7901
rect 3030 7842 3076 7854
rect 3030 7766 3036 7842
rect 3070 7766 3076 7842
rect 3030 7754 3076 7766
rect 3488 7842 3534 7854
rect 3488 7766 3494 7842
rect 3528 7766 3534 7842
rect 3488 7754 3534 7766
rect 3730 7842 3776 7854
rect 3730 7766 3736 7842
rect 3770 7766 3776 7842
rect 3730 7754 3776 7766
rect 4188 7842 4234 7854
rect 4188 7766 4194 7842
rect 4228 7766 4234 7842
rect 4188 7754 4234 7766
rect 59 7595 2765 7695
rect 3086 7707 3478 7713
rect 3086 7673 3098 7707
rect 3466 7673 3478 7707
rect 3086 7667 3478 7673
rect 3786 7707 4178 7713
rect 3786 7673 3798 7707
rect 4166 7673 4178 7707
rect 3786 7667 4178 7673
rect -347 7580 2765 7595
rect -347 7575 1167 7580
rect -347 7573 1105 7575
rect -347 7545 116 7573
rect 4766 7246 4854 9676
rect 5270 7246 5354 9676
rect 5810 9753 5852 9961
rect 5930 9945 7030 9951
rect 5930 9911 5942 9945
rect 7018 9911 7030 9945
rect 5930 9905 7030 9911
rect 5930 9803 7030 9809
rect 5930 9769 5942 9803
rect 7018 9769 7030 9803
rect 5930 9763 7030 9769
rect 7108 9755 7150 9961
rect 7376 9899 8476 9905
rect 7376 9865 7388 9899
rect 8464 9865 8476 9899
rect 7376 9859 8476 9865
rect 8714 9858 8749 9973
rect 8976 9956 8982 10084
rect 9016 9956 9022 10084
rect 8976 9944 9022 9956
rect 9304 10084 9350 10096
rect 9304 9956 9310 10084
rect 9344 9956 9350 10084
rect 9304 9944 9350 9956
rect 9667 10084 9713 10096
rect 9667 9956 9673 10084
rect 9707 9956 9713 10084
rect 9667 9944 9713 9956
rect 9995 10084 10041 10096
rect 9995 9956 10001 10084
rect 10035 9956 10041 10084
rect 10215 10081 10234 10164
rect 10269 10081 10287 10164
rect 10215 10065 10287 10081
rect 10385 10223 11737 10267
rect 10385 10131 10433 10223
rect 10511 10181 11611 10187
rect 10511 10147 10523 10181
rect 11599 10147 11611 10181
rect 10511 10141 11611 10147
rect 11689 10131 11737 10223
rect 10385 10119 10479 10131
rect 10385 10071 10439 10119
rect 10473 10071 10479 10119
rect 10385 10059 10479 10071
rect 11643 10119 11737 10131
rect 11643 10071 11649 10119
rect 11683 10071 11737 10119
rect 11643 10059 11737 10071
rect 11867 10461 11955 10473
rect 11867 10333 11915 10461
rect 11949 10333 11955 10461
rect 11867 10321 11955 10333
rect 13119 10461 13207 10473
rect 13119 10333 13125 10461
rect 13159 10333 13207 10461
rect 13119 10321 13207 10333
rect 11867 10113 11909 10321
rect 11987 10305 13087 10311
rect 11987 10271 11999 10305
rect 13075 10271 13087 10305
rect 11987 10265 13087 10271
rect 11987 10163 13087 10169
rect 11987 10129 11999 10163
rect 13075 10129 13087 10163
rect 11987 10123 13087 10129
rect 13165 10113 13207 10321
rect 11867 10101 11955 10113
rect 10511 10043 11611 10049
rect 10511 10014 10523 10043
rect 9995 9944 10041 9956
rect 10268 10009 10523 10014
rect 11599 10009 11611 10043
rect 10268 10003 11611 10009
rect 10268 9973 10768 10003
rect 11867 9973 11915 10101
rect 11949 9973 11955 10101
rect 9063 9928 9263 9934
rect 9063 9894 9075 9928
rect 9251 9894 9263 9928
rect 9063 9888 9263 9894
rect 9754 9928 9954 9934
rect 9754 9894 9766 9928
rect 9942 9894 9954 9928
rect 9754 9888 9954 9894
rect 9126 9858 9196 9888
rect 7256 9837 7344 9849
rect 7256 9755 7304 9837
rect 7108 9753 7304 9755
rect 5810 9741 5898 9753
rect 5810 9613 5858 9741
rect 5892 9613 5898 9741
rect 5810 9601 5898 9613
rect 7062 9741 7304 9753
rect 7062 9613 7068 9741
rect 7102 9693 7304 9741
rect 7102 9645 7150 9693
rect 7256 9669 7304 9693
rect 7338 9669 7344 9837
rect 7256 9657 7344 9669
rect 8508 9837 8596 9849
rect 8508 9669 8514 9837
rect 8548 9669 8596 9837
rect 8714 9774 9196 9858
rect 9821 9858 9891 9888
rect 10268 9858 10303 9973
rect 11867 9961 11955 9973
rect 13119 10101 13207 10113
rect 13119 9973 13125 10101
rect 13159 9973 13207 10101
rect 13119 9961 13207 9973
rect 10541 9899 11641 9905
rect 10541 9865 10553 9899
rect 11629 9865 11641 9899
rect 10541 9859 11641 9865
rect 9126 9706 9196 9774
rect 9271 9831 9376 9853
rect 9271 9763 9291 9831
rect 9354 9763 9376 9831
rect 9271 9746 9376 9763
rect 9641 9831 9746 9853
rect 9641 9763 9663 9831
rect 9726 9763 9746 9831
rect 9641 9746 9746 9763
rect 9821 9774 10303 9858
rect 10421 9837 10509 9849
rect 9821 9706 9891 9774
rect 8508 9657 8596 9669
rect 9063 9700 9263 9706
rect 9063 9666 9075 9700
rect 9251 9666 9263 9700
rect 9063 9660 9263 9666
rect 9754 9700 9954 9706
rect 9754 9666 9766 9700
rect 9942 9666 9954 9700
rect 9754 9660 9954 9666
rect 10421 9669 10469 9837
rect 10503 9669 10509 9837
rect 7102 9613 7152 9645
rect 7062 9601 7152 9613
rect 5810 9393 5852 9601
rect 5930 9585 7030 9591
rect 5930 9551 5942 9585
rect 7018 9551 7030 9585
rect 5930 9545 7030 9551
rect 5930 9443 7030 9449
rect 5930 9409 5942 9443
rect 7018 9409 7030 9443
rect 5930 9403 7030 9409
rect 7108 9425 7152 9601
rect 7256 9563 7298 9657
rect 7376 9641 8476 9647
rect 7376 9607 7388 9641
rect 8464 9607 8476 9641
rect 7376 9601 8476 9607
rect 8554 9563 8596 9657
rect 10421 9657 10509 9669
rect 11673 9837 11761 9849
rect 11673 9669 11679 9837
rect 11713 9755 11761 9837
rect 11867 9755 11909 9961
rect 11987 9945 13087 9951
rect 11987 9911 11999 9945
rect 13075 9911 13087 9945
rect 11987 9905 13087 9911
rect 11987 9803 13087 9809
rect 11987 9769 11999 9803
rect 13075 9769 13087 9803
rect 11987 9763 13087 9769
rect 11713 9753 11909 9755
rect 13165 9753 13207 9961
rect 11713 9741 11955 9753
rect 11713 9693 11915 9741
rect 11713 9669 11761 9693
rect 11673 9657 11761 9669
rect 7256 9525 8596 9563
rect 7256 9425 7298 9525
rect 7376 9475 8476 9481
rect 7376 9441 7388 9475
rect 8464 9441 8476 9475
rect 7376 9435 8476 9441
rect 8554 9432 8596 9525
rect 8976 9638 9022 9650
rect 8976 9432 8982 9638
rect 8554 9425 8982 9432
rect 7108 9393 7150 9425
rect 5810 9381 5898 9393
rect 5810 9253 5858 9381
rect 5892 9253 5898 9381
rect 5810 9241 5898 9253
rect 7062 9381 7150 9393
rect 7062 9253 7068 9381
rect 7102 9371 7150 9381
rect 7256 9413 7344 9425
rect 7256 9371 7304 9413
rect 7102 9309 7304 9371
rect 7102 9253 7150 9309
rect 7062 9241 7150 9253
rect 7256 9245 7304 9309
rect 7338 9245 7344 9413
rect 7256 9233 7344 9245
rect 8508 9413 8982 9425
rect 8508 9245 8514 9413
rect 8548 9299 8982 9413
rect 8548 9245 8596 9299
rect 8976 9270 8982 9299
rect 9016 9270 9022 9638
rect 8976 9258 9022 9270
rect 9304 9638 9350 9650
rect 9304 9270 9310 9638
rect 9344 9270 9350 9638
rect 9304 9258 9350 9270
rect 9667 9638 9713 9650
rect 9667 9270 9673 9638
rect 9707 9270 9713 9638
rect 9667 9258 9713 9270
rect 9995 9638 10041 9650
rect 9995 9270 10001 9638
rect 10035 9432 10041 9638
rect 10421 9563 10463 9657
rect 10541 9641 11641 9647
rect 10541 9607 10553 9641
rect 11629 9607 11641 9641
rect 10541 9601 11641 9607
rect 11719 9563 11761 9657
rect 11867 9645 11915 9693
rect 10421 9525 11761 9563
rect 10421 9432 10463 9525
rect 10541 9475 11641 9481
rect 10541 9441 10553 9475
rect 11629 9441 11641 9475
rect 10541 9435 11641 9441
rect 10035 9425 10463 9432
rect 11719 9425 11761 9525
rect 11865 9613 11915 9645
rect 11949 9613 11955 9741
rect 11865 9601 11955 9613
rect 13119 9741 13207 9753
rect 13119 9613 13125 9741
rect 13159 9613 13207 9741
rect 13119 9601 13207 9613
rect 11865 9425 11909 9601
rect 11987 9585 13087 9591
rect 11987 9551 11999 9585
rect 13075 9551 13087 9585
rect 11987 9545 13087 9551
rect 10035 9413 10509 9425
rect 10035 9299 10469 9413
rect 10035 9270 10041 9299
rect 9995 9258 10041 9270
rect 8508 9233 8596 9245
rect 9063 9242 9263 9248
rect 5930 9225 7030 9231
rect 5930 9191 5942 9225
rect 7018 9191 7030 9225
rect 5930 9185 7030 9191
rect 7376 9217 8476 9223
rect 7376 9183 7388 9217
rect 8464 9183 8476 9217
rect 9063 9208 9075 9242
rect 9251 9208 9263 9242
rect 9063 9202 9263 9208
rect 9754 9242 9954 9248
rect 9754 9208 9766 9242
rect 9942 9208 9954 9242
rect 10421 9245 10469 9299
rect 10503 9245 10509 9413
rect 10421 9233 10509 9245
rect 11673 9413 11761 9425
rect 11673 9245 11679 9413
rect 11713 9371 11761 9413
rect 11867 9393 11909 9425
rect 11987 9443 13087 9449
rect 11987 9409 11999 9443
rect 13075 9409 13087 9443
rect 11987 9403 13087 9409
rect 13165 9393 13207 9601
rect 11867 9381 11955 9393
rect 11867 9371 11915 9381
rect 11713 9309 11915 9371
rect 11713 9245 11761 9309
rect 11673 9233 11761 9245
rect 11867 9253 11915 9309
rect 11949 9253 11955 9381
rect 11867 9241 11955 9253
rect 13119 9381 13207 9393
rect 13119 9253 13125 9381
rect 13159 9253 13207 9381
rect 13119 9241 13207 9253
rect 11987 9225 13087 9231
rect 9754 9202 9954 9208
rect 10541 9217 11641 9223
rect 7376 9177 8476 9183
rect 10541 9183 10553 9217
rect 11629 9183 11641 9217
rect 11987 9191 11999 9225
rect 13075 9191 13087 9225
rect 11987 9185 13087 9191
rect 10541 9177 11641 9183
rect 8388 9060 8672 9061
rect 10345 9060 10629 9061
rect 8388 9043 9189 9060
rect 8388 8974 8416 9043
rect 8643 8974 9189 9043
rect 8388 8971 9189 8974
rect 8388 8961 8672 8971
rect 7125 8897 7330 8939
rect 6450 8863 8801 8897
rect 9130 8894 9189 8971
rect 9828 9043 10629 9060
rect 9828 8974 10374 9043
rect 10601 8974 10629 9043
rect 9828 8971 10629 8974
rect 9828 8894 9887 8971
rect 10345 8961 10629 8971
rect 11687 8897 11892 8939
rect 5930 8861 8801 8863
rect 5930 8857 7030 8861
rect 5930 8823 5942 8857
rect 7018 8823 7030 8857
rect 5930 8817 7030 8823
rect 7280 8857 8801 8861
rect 5810 8795 5898 8807
rect 5810 8667 5858 8795
rect 5892 8667 5898 8795
rect 5810 8655 5898 8667
rect 7062 8795 7150 8807
rect 7062 8667 7068 8795
rect 7102 8667 7150 8795
rect 7062 8655 7150 8667
rect 5810 8447 5852 8655
rect 5930 8639 7030 8645
rect 5930 8605 5942 8639
rect 7018 8605 7030 8639
rect 5930 8599 7030 8605
rect 5930 8497 7030 8503
rect 5930 8463 5942 8497
rect 7018 8463 7030 8497
rect 5930 8457 7030 8463
rect 7108 8447 7150 8655
rect 5810 8435 5898 8447
rect 5810 8307 5858 8435
rect 5892 8307 5898 8435
rect 5810 8295 5898 8307
rect 7062 8435 7150 8447
rect 7062 8307 7068 8435
rect 7102 8307 7150 8435
rect 7280 8763 7328 8857
rect 8733 8828 8801 8857
rect 9063 8888 9263 8894
rect 9063 8854 9075 8888
rect 9251 8854 9263 8888
rect 9063 8848 9263 8854
rect 9754 8888 9954 8894
rect 9754 8854 9766 8888
rect 9942 8854 9954 8888
rect 9754 8848 9954 8854
rect 10216 8863 12567 8897
rect 10216 8861 13087 8863
rect 10216 8857 11737 8861
rect 8976 8828 9022 8838
rect 8733 8826 9022 8828
rect 7406 8813 8506 8819
rect 7406 8779 7418 8813
rect 8494 8779 8506 8813
rect 7406 8773 8506 8779
rect 8733 8768 8982 8826
rect 8733 8767 8801 8768
rect 7280 8751 7374 8763
rect 7280 8703 7334 8751
rect 7368 8703 7374 8751
rect 7280 8691 7374 8703
rect 8538 8751 8632 8763
rect 8538 8703 8544 8751
rect 8578 8703 8632 8751
rect 8538 8691 8632 8703
rect 7280 8601 7328 8691
rect 7406 8675 8506 8681
rect 7406 8641 7418 8675
rect 8494 8641 8506 8675
rect 7406 8635 8506 8641
rect 8584 8601 8632 8691
rect 8976 8698 8982 8768
rect 9016 8698 9022 8826
rect 8976 8686 9022 8698
rect 9304 8826 9350 8838
rect 9304 8698 9310 8826
rect 9344 8698 9350 8826
rect 9304 8686 9350 8698
rect 9667 8826 9713 8838
rect 9667 8698 9673 8826
rect 9707 8698 9713 8826
rect 9667 8686 9713 8698
rect 9995 8828 10041 8838
rect 10216 8828 10284 8857
rect 9995 8826 10284 8828
rect 9995 8698 10001 8826
rect 10035 8768 10284 8826
rect 10511 8813 11611 8819
rect 10511 8779 10523 8813
rect 11599 8779 11611 8813
rect 10511 8773 11611 8779
rect 10035 8698 10041 8768
rect 10216 8767 10284 8768
rect 11689 8763 11737 8857
rect 11987 8857 13087 8861
rect 11987 8823 11999 8857
rect 13075 8823 13087 8857
rect 11987 8817 13087 8823
rect 9995 8686 10041 8698
rect 10385 8751 10479 8763
rect 10385 8703 10439 8751
rect 10473 8703 10479 8751
rect 10385 8691 10479 8703
rect 11643 8751 11737 8763
rect 11643 8703 11649 8751
rect 11683 8703 11737 8751
rect 11643 8691 11737 8703
rect 9063 8670 9263 8676
rect 9063 8636 9075 8670
rect 9251 8636 9263 8670
rect 9063 8630 9263 8636
rect 9754 8670 9954 8676
rect 9754 8636 9766 8670
rect 9942 8636 9954 8670
rect 9754 8630 9954 8636
rect 7280 8557 8632 8601
rect 9143 8575 9187 8630
rect 7280 8465 7328 8557
rect 7406 8515 8506 8521
rect 7406 8481 7418 8515
rect 8494 8481 8506 8515
rect 7406 8475 8506 8481
rect 8584 8465 8632 8557
rect 7280 8453 7374 8465
rect 7280 8405 7334 8453
rect 7368 8405 7374 8453
rect 7280 8393 7374 8405
rect 8538 8453 8632 8465
rect 8538 8405 8544 8453
rect 8578 8405 8632 8453
rect 8538 8393 8632 8405
rect 8730 8530 9187 8575
rect 9249 8582 9436 8600
rect 9249 8530 9274 8582
rect 9372 8530 9436 8582
rect 8730 8498 8802 8530
rect 9249 8515 9436 8530
rect 9581 8582 9768 8600
rect 9581 8530 9645 8582
rect 9743 8530 9768 8582
rect 9830 8575 9874 8630
rect 10385 8601 10433 8691
rect 10511 8675 11611 8681
rect 10511 8641 10523 8675
rect 11599 8641 11611 8675
rect 10511 8635 11611 8641
rect 11689 8601 11737 8691
rect 9830 8530 10287 8575
rect 9581 8515 9768 8530
rect 8730 8415 8748 8498
rect 8783 8415 8802 8498
rect 10215 8498 10287 8530
rect 9063 8480 9263 8486
rect 9063 8446 9075 8480
rect 9251 8446 9263 8480
rect 9063 8440 9263 8446
rect 9754 8480 9954 8486
rect 9754 8446 9766 8480
rect 9942 8446 9954 8480
rect 9754 8440 9954 8446
rect 8730 8399 8802 8415
rect 8976 8418 9022 8430
rect 7406 8377 8506 8383
rect 7406 8343 7418 8377
rect 8494 8348 8506 8377
rect 8494 8343 8749 8348
rect 7406 8337 8749 8343
rect 8249 8307 8749 8337
rect 7062 8295 7150 8307
rect 5810 8087 5852 8295
rect 5930 8279 7030 8285
rect 5930 8245 5942 8279
rect 7018 8245 7030 8279
rect 5930 8239 7030 8245
rect 5930 8137 7030 8143
rect 5930 8103 5942 8137
rect 7018 8103 7030 8137
rect 5930 8097 7030 8103
rect 7108 8089 7150 8295
rect 7376 8233 8476 8239
rect 7376 8199 7388 8233
rect 8464 8199 8476 8233
rect 7376 8193 8476 8199
rect 8714 8192 8749 8307
rect 8976 8290 8982 8418
rect 9016 8290 9022 8418
rect 8976 8278 9022 8290
rect 9304 8418 9350 8430
rect 9304 8290 9310 8418
rect 9344 8290 9350 8418
rect 9304 8278 9350 8290
rect 9667 8418 9713 8430
rect 9667 8290 9673 8418
rect 9707 8290 9713 8418
rect 9667 8278 9713 8290
rect 9995 8418 10041 8430
rect 9995 8290 10001 8418
rect 10035 8290 10041 8418
rect 10215 8415 10234 8498
rect 10269 8415 10287 8498
rect 10215 8399 10287 8415
rect 10385 8557 11737 8601
rect 10385 8465 10433 8557
rect 10511 8515 11611 8521
rect 10511 8481 10523 8515
rect 11599 8481 11611 8515
rect 10511 8475 11611 8481
rect 11689 8465 11737 8557
rect 10385 8453 10479 8465
rect 10385 8405 10439 8453
rect 10473 8405 10479 8453
rect 10385 8393 10479 8405
rect 11643 8453 11737 8465
rect 11643 8405 11649 8453
rect 11683 8405 11737 8453
rect 11643 8393 11737 8405
rect 11867 8795 11955 8807
rect 11867 8667 11915 8795
rect 11949 8667 11955 8795
rect 11867 8655 11955 8667
rect 13119 8795 13207 8807
rect 13119 8667 13125 8795
rect 13159 8667 13207 8795
rect 13119 8655 13207 8667
rect 11867 8447 11909 8655
rect 11987 8639 13087 8645
rect 11987 8605 11999 8639
rect 13075 8605 13087 8639
rect 11987 8599 13087 8605
rect 11987 8497 13087 8503
rect 11987 8463 11999 8497
rect 13075 8463 13087 8497
rect 11987 8457 13087 8463
rect 13165 8447 13207 8655
rect 11867 8435 11955 8447
rect 10511 8377 11611 8383
rect 10511 8348 10523 8377
rect 9995 8278 10041 8290
rect 10268 8343 10523 8348
rect 11599 8343 11611 8377
rect 10268 8337 11611 8343
rect 10268 8307 10768 8337
rect 11867 8307 11915 8435
rect 11949 8307 11955 8435
rect 9063 8262 9263 8268
rect 9063 8228 9075 8262
rect 9251 8228 9263 8262
rect 9063 8222 9263 8228
rect 9754 8262 9954 8268
rect 9754 8228 9766 8262
rect 9942 8228 9954 8262
rect 9754 8222 9954 8228
rect 9126 8192 9196 8222
rect 7256 8171 7344 8183
rect 7256 8089 7304 8171
rect 7108 8087 7304 8089
rect 5810 8075 5898 8087
rect 5810 7947 5858 8075
rect 5892 7947 5898 8075
rect 5810 7935 5898 7947
rect 7062 8075 7304 8087
rect 7062 7947 7068 8075
rect 7102 8027 7304 8075
rect 7102 7979 7150 8027
rect 7256 8003 7304 8027
rect 7338 8003 7344 8171
rect 7256 7991 7344 8003
rect 8508 8171 8596 8183
rect 8508 8003 8514 8171
rect 8548 8003 8596 8171
rect 8714 8108 9196 8192
rect 9821 8192 9891 8222
rect 10268 8192 10303 8307
rect 11867 8295 11955 8307
rect 13119 8435 13207 8447
rect 13119 8307 13125 8435
rect 13159 8307 13207 8435
rect 13119 8295 13207 8307
rect 10541 8233 11641 8239
rect 10541 8199 10553 8233
rect 11629 8199 11641 8233
rect 10541 8193 11641 8199
rect 9126 8040 9196 8108
rect 9271 8165 9376 8187
rect 9271 8097 9291 8165
rect 9354 8097 9376 8165
rect 9271 8080 9376 8097
rect 9641 8165 9746 8187
rect 9641 8097 9663 8165
rect 9726 8097 9746 8165
rect 9641 8080 9746 8097
rect 9821 8108 10303 8192
rect 10421 8171 10509 8183
rect 9821 8040 9891 8108
rect 8508 7991 8596 8003
rect 9063 8034 9263 8040
rect 9063 8000 9075 8034
rect 9251 8000 9263 8034
rect 9063 7994 9263 8000
rect 9754 8034 9954 8040
rect 9754 8000 9766 8034
rect 9942 8000 9954 8034
rect 9754 7994 9954 8000
rect 10421 8003 10469 8171
rect 10503 8003 10509 8171
rect 7102 7947 7152 7979
rect 7062 7935 7152 7947
rect 5810 7727 5852 7935
rect 5930 7919 7030 7925
rect 5930 7885 5942 7919
rect 7018 7885 7030 7919
rect 5930 7879 7030 7885
rect 5930 7777 7030 7783
rect 5930 7743 5942 7777
rect 7018 7743 7030 7777
rect 5930 7737 7030 7743
rect 7108 7759 7152 7935
rect 7256 7897 7298 7991
rect 7376 7975 8476 7981
rect 7376 7941 7388 7975
rect 8464 7941 8476 7975
rect 7376 7935 8476 7941
rect 8554 7897 8596 7991
rect 10421 7991 10509 8003
rect 11673 8171 11761 8183
rect 11673 8003 11679 8171
rect 11713 8089 11761 8171
rect 11867 8089 11909 8295
rect 11987 8279 13087 8285
rect 11987 8245 11999 8279
rect 13075 8245 13087 8279
rect 11987 8239 13087 8245
rect 11987 8137 13087 8143
rect 11987 8103 11999 8137
rect 13075 8103 13087 8137
rect 11987 8097 13087 8103
rect 11713 8087 11909 8089
rect 13165 8087 13207 8295
rect 11713 8075 11955 8087
rect 11713 8027 11915 8075
rect 11713 8003 11761 8027
rect 11673 7991 11761 8003
rect 7256 7859 8596 7897
rect 7256 7759 7298 7859
rect 7376 7809 8476 7815
rect 7376 7775 7388 7809
rect 8464 7775 8476 7809
rect 7376 7769 8476 7775
rect 8554 7766 8596 7859
rect 8976 7972 9022 7984
rect 8976 7766 8982 7972
rect 8554 7759 8982 7766
rect 7108 7727 7150 7759
rect 5810 7715 5898 7727
rect 5810 7587 5858 7715
rect 5892 7587 5898 7715
rect 5810 7575 5898 7587
rect 7062 7715 7150 7727
rect 7062 7587 7068 7715
rect 7102 7705 7150 7715
rect 7256 7747 7344 7759
rect 7256 7705 7304 7747
rect 7102 7643 7304 7705
rect 7102 7587 7150 7643
rect 7062 7575 7150 7587
rect 7256 7579 7304 7643
rect 7338 7579 7344 7747
rect 7256 7567 7344 7579
rect 8508 7747 8982 7759
rect 8508 7579 8514 7747
rect 8548 7633 8982 7747
rect 8548 7579 8596 7633
rect 8976 7604 8982 7633
rect 9016 7604 9022 7972
rect 8976 7592 9022 7604
rect 9304 7972 9350 7984
rect 9304 7604 9310 7972
rect 9344 7604 9350 7972
rect 9304 7592 9350 7604
rect 9667 7972 9713 7984
rect 9667 7604 9673 7972
rect 9707 7604 9713 7972
rect 9667 7592 9713 7604
rect 9995 7972 10041 7984
rect 9995 7604 10001 7972
rect 10035 7766 10041 7972
rect 10421 7897 10463 7991
rect 10541 7975 11641 7981
rect 10541 7941 10553 7975
rect 11629 7941 11641 7975
rect 10541 7935 11641 7941
rect 11719 7897 11761 7991
rect 11867 7979 11915 8027
rect 10421 7859 11761 7897
rect 10421 7766 10463 7859
rect 10541 7809 11641 7815
rect 10541 7775 10553 7809
rect 11629 7775 11641 7809
rect 10541 7769 11641 7775
rect 10035 7759 10463 7766
rect 11719 7759 11761 7859
rect 11865 7947 11915 7979
rect 11949 7947 11955 8075
rect 11865 7935 11955 7947
rect 13119 8075 13207 8087
rect 13119 7947 13125 8075
rect 13159 7947 13207 8075
rect 13119 7935 13207 7947
rect 11865 7759 11909 7935
rect 11987 7919 13087 7925
rect 11987 7885 11999 7919
rect 13075 7885 13087 7919
rect 11987 7879 13087 7885
rect 10035 7747 10509 7759
rect 10035 7633 10469 7747
rect 10035 7604 10041 7633
rect 9995 7592 10041 7604
rect 8508 7567 8596 7579
rect 9063 7576 9263 7582
rect 5930 7559 7030 7565
rect 5930 7525 5942 7559
rect 7018 7525 7030 7559
rect 5930 7519 7030 7525
rect 7376 7551 8476 7557
rect 7376 7517 7388 7551
rect 8464 7517 8476 7551
rect 9063 7542 9075 7576
rect 9251 7542 9263 7576
rect 9063 7536 9263 7542
rect 9754 7576 9954 7582
rect 9754 7542 9766 7576
rect 9942 7542 9954 7576
rect 10421 7579 10469 7633
rect 10503 7579 10509 7747
rect 10421 7567 10509 7579
rect 11673 7747 11761 7759
rect 11673 7579 11679 7747
rect 11713 7705 11761 7747
rect 11867 7727 11909 7759
rect 11987 7777 13087 7783
rect 11987 7743 11999 7777
rect 13075 7743 13087 7777
rect 11987 7737 13087 7743
rect 13165 7727 13207 7935
rect 11867 7715 11955 7727
rect 11867 7705 11915 7715
rect 11713 7643 11915 7705
rect 11713 7579 11761 7643
rect 11673 7567 11761 7579
rect 11867 7587 11915 7643
rect 11949 7587 11955 7715
rect 11867 7575 11955 7587
rect 13119 7715 13207 7727
rect 13119 7587 13125 7715
rect 13159 7587 13207 7715
rect 13119 7575 13207 7587
rect 11987 7559 13087 7565
rect 9754 7536 9954 7542
rect 10541 7551 11641 7557
rect 7376 7511 8476 7517
rect 10541 7517 10553 7551
rect 11629 7517 11641 7551
rect 11987 7525 11999 7559
rect 13075 7525 13087 7559
rect 11987 7519 13087 7525
rect 10541 7511 11641 7517
rect 4766 7166 5354 7246
rect 4766 6140 5352 7166
rect 13599 6140 14090 13882
rect 17989 13660 18511 13886
rect 17988 13538 18511 13660
rect 14982 13502 15160 13508
rect 14982 13468 14994 13502
rect 15148 13468 15160 13502
rect 14982 13462 15160 13468
rect 15482 13502 15660 13508
rect 15482 13468 15494 13502
rect 15648 13468 15660 13502
rect 15482 13462 15660 13468
rect 15982 13502 16160 13508
rect 15982 13468 15994 13502
rect 16148 13468 16160 13502
rect 15982 13462 16160 13468
rect 16482 13502 16660 13508
rect 16482 13468 16494 13502
rect 16648 13468 16660 13502
rect 16482 13462 16660 13468
rect 16982 13502 17160 13508
rect 16982 13468 16994 13502
rect 17148 13468 17160 13502
rect 16982 13462 17160 13468
rect 17482 13502 17660 13508
rect 17482 13468 17494 13502
rect 17648 13468 17660 13502
rect 17482 13462 17660 13468
rect 14895 13440 14941 13452
rect 14895 12694 14901 13440
rect 14935 12694 14941 13440
rect 14895 12682 14941 12694
rect 15201 13440 15247 13452
rect 15201 12694 15207 13440
rect 15241 12694 15247 13440
rect 15201 12682 15247 12694
rect 15395 13440 15441 13452
rect 15395 12694 15401 13440
rect 15435 12694 15441 13440
rect 15395 12682 15441 12694
rect 15701 13440 15747 13452
rect 15701 12694 15707 13440
rect 15741 13132 15747 13440
rect 15895 13440 15941 13452
rect 15895 13132 15901 13440
rect 15741 12998 15901 13132
rect 15741 12694 15747 12998
rect 15701 12682 15747 12694
rect 15895 12694 15901 12998
rect 15935 12694 15941 13440
rect 15895 12682 15941 12694
rect 16201 13440 16247 13452
rect 16201 12694 16207 13440
rect 16241 13132 16247 13440
rect 16395 13440 16441 13452
rect 16395 13132 16401 13440
rect 16241 12998 16401 13132
rect 16241 12869 16247 12998
rect 16395 12869 16401 12998
rect 16241 12815 16401 12869
rect 16241 12694 16258 12815
rect 16201 12682 16258 12694
rect 16160 12672 16258 12682
rect 14982 12666 15160 12672
rect 14982 12632 14994 12666
rect 15148 12632 15160 12666
rect 14982 12626 15160 12632
rect 15482 12666 15660 12672
rect 15482 12632 15494 12666
rect 15648 12632 15660 12666
rect 15482 12626 15660 12632
rect 15982 12666 16258 12672
rect 15982 12632 15994 12666
rect 16148 12664 16258 12666
rect 16384 12694 16401 12815
rect 16435 12694 16441 13440
rect 16384 12682 16441 12694
rect 16701 13440 16747 13452
rect 16701 12694 16707 13440
rect 16741 13132 16747 13440
rect 16895 13440 16941 13452
rect 16895 13132 16901 13440
rect 16741 12998 16901 13132
rect 16741 12694 16747 12998
rect 16701 12682 16747 12694
rect 16895 12694 16901 12998
rect 16935 12694 16941 13440
rect 16895 12682 16941 12694
rect 17201 13440 17247 13452
rect 17201 12694 17207 13440
rect 17241 12694 17247 13440
rect 17201 12682 17247 12694
rect 17395 13440 17441 13452
rect 17395 12694 17401 13440
rect 17435 12694 17441 13440
rect 17395 12682 17441 12694
rect 17701 13440 17747 13452
rect 17701 12694 17707 13440
rect 17741 12694 17747 13440
rect 17701 12682 17747 12694
rect 16384 12672 16482 12682
rect 16384 12666 16660 12672
rect 16384 12664 16494 12666
rect 16148 12632 16494 12664
rect 16648 12632 16660 12666
rect 15982 12626 16660 12632
rect 16982 12666 17160 12672
rect 16982 12632 16994 12666
rect 17148 12632 17160 12666
rect 16982 12626 17160 12632
rect 17482 12666 17660 12672
rect 17482 12632 17494 12666
rect 17648 12632 17660 12666
rect 17482 12626 17660 12632
rect 15544 12559 15604 12626
rect 17044 12559 17104 12626
rect 14899 12532 15418 12555
rect 14899 12442 14975 12532
rect 15349 12442 15418 12532
rect 15544 12509 17104 12559
rect 14899 12422 15418 12442
rect 14340 12225 14787 12298
rect 14340 12043 14431 12225
rect 14693 12043 14787 12225
rect 14340 11971 14787 12043
rect 14355 11674 14462 11971
rect 14552 11768 15198 11814
rect 14552 11752 15078 11768
rect 14552 11746 14830 11752
rect 14552 11712 14564 11746
rect 14818 11712 14830 11746
rect 14552 11706 14830 11712
rect 14355 11662 14542 11674
rect 14355 10648 14502 11662
rect 14536 10648 14542 11662
rect 14355 10636 14542 10648
rect 14840 11662 14886 11674
rect 14840 10648 14846 11662
rect 14880 11566 14886 11662
rect 14880 11536 14952 11566
rect 14924 10673 14952 11536
rect 14880 10648 14952 10673
rect 14840 10636 14952 10648
rect 15042 11092 15078 11752
rect 15159 11092 15198 11768
rect 15042 11050 15198 11092
rect 14355 10418 14496 10636
rect 14552 10598 14830 10604
rect 14552 10564 14564 10598
rect 14818 10564 14830 10598
rect 14552 10558 14830 10564
rect 15042 10558 15094 11050
rect 14552 10496 15094 10558
rect 14552 10490 14830 10496
rect 14552 10456 14564 10490
rect 14818 10456 14830 10490
rect 14552 10450 14830 10456
rect 14355 10406 14542 10418
rect 14355 10331 14502 10406
rect 14446 9392 14502 10331
rect 14536 9392 14542 10406
rect 14446 9380 14542 9392
rect 14840 10406 14952 10418
rect 14840 9392 14846 10406
rect 14880 10382 14952 10406
rect 14919 9519 14952 10382
rect 14880 9488 14952 9519
rect 14880 9392 14886 9488
rect 14840 9380 14886 9392
rect 14552 9342 14830 9348
rect 14552 9308 14564 9342
rect 14818 9308 14830 9342
rect 14552 9302 14830 9308
rect 15042 9302 15094 10496
rect 14552 9240 15094 9302
rect 15320 9043 15415 12422
rect 16532 12382 16664 12509
rect 16532 12264 16562 12382
rect 16633 12264 16664 12382
rect 16532 12226 16664 12264
rect 17988 12101 18062 13538
rect 18236 13054 18511 13538
rect 18236 12101 18317 13054
rect 17988 11988 18317 12101
rect 16722 11549 18207 11583
rect 16722 11266 16750 11549
rect 16829 11536 18207 11549
rect 16829 11289 16857 11536
rect 17086 11347 18120 11353
rect 17086 11313 17098 11347
rect 18108 11313 18120 11347
rect 17086 11307 18120 11313
rect 16999 11289 17045 11297
rect 16829 11285 17045 11289
rect 16829 11266 17005 11285
rect 16722 11243 17005 11266
rect 17039 11243 17045 11285
rect 16722 11233 17045 11243
rect 16999 11231 17045 11233
rect 18161 11285 18207 11536
rect 18161 11243 18167 11285
rect 18201 11243 18207 11285
rect 18161 11231 18207 11243
rect 17086 11215 18120 11221
rect 17086 11181 17098 11215
rect 18108 11181 18120 11215
rect 17086 11175 18120 11181
rect 17530 10988 17652 11175
rect 17058 10984 17654 10988
rect 17851 10984 18686 10994
rect 17058 10942 18686 10984
rect 17058 10640 17124 10942
rect 17596 10764 18686 10942
rect 17596 10667 17654 10764
rect 17596 10640 17709 10667
rect 17058 10602 17709 10640
rect 17058 10592 17513 10602
rect 17481 10353 17513 10592
rect 16815 10323 17513 10353
rect 17670 10353 17709 10602
rect 17851 10566 18686 10764
rect 18067 10565 18686 10566
rect 17670 10323 18243 10353
rect 16815 10286 18243 10323
rect 16815 9753 16902 10286
rect 17029 10280 18243 10286
rect 17029 10246 17041 10280
rect 18231 10246 18243 10280
rect 17029 10240 18243 10246
rect 16942 10218 16988 10230
rect 16942 9996 16948 10218
rect 16982 9996 16988 10218
rect 16942 9984 16988 9996
rect 18284 10218 18330 10230
rect 18284 9996 18290 10218
rect 18324 10212 18330 10218
rect 18401 10212 18782 10214
rect 18324 10012 18782 10212
rect 18324 9996 18330 10012
rect 18401 10009 18782 10012
rect 18284 9984 18330 9996
rect 17029 9968 18243 9974
rect 17029 9934 17041 9968
rect 18231 9934 18243 9968
rect 17029 9928 18243 9934
rect 17029 9861 18463 9928
rect 16815 9686 18243 9753
rect 17029 9680 18243 9686
rect 17029 9646 17041 9680
rect 18231 9646 18243 9680
rect 17029 9640 18243 9646
rect 16942 9618 16988 9630
rect 16942 9396 16948 9618
rect 16982 9396 16988 9618
rect 16942 9384 16988 9396
rect 18284 9618 18330 9630
rect 18284 9396 18290 9618
rect 18324 9396 18330 9618
rect 18284 9384 18330 9396
rect 17029 9368 18243 9374
rect 17029 9334 17041 9368
rect 18231 9334 18243 9368
rect 17029 9328 18243 9334
rect 18376 9328 18463 9861
rect 17029 9326 18463 9328
rect 17027 9283 18463 9326
rect 17027 9153 17058 9283
rect 17230 9261 18463 9283
rect 17230 9153 17271 9261
rect 17027 9133 17271 9153
rect 15106 8990 17670 9043
rect 14526 8670 14650 8676
rect 14526 8636 14538 8670
rect 14638 8636 14650 8670
rect 14526 8630 14650 8636
rect 14926 8670 15050 8676
rect 14926 8636 14938 8670
rect 15038 8636 15050 8670
rect 14926 8630 15050 8636
rect 15106 8598 15161 8990
rect 15506 8879 17270 8920
rect 15506 8792 15580 8879
rect 15879 8872 16890 8879
rect 15879 8792 15961 8872
rect 15506 8750 15961 8792
rect 15326 8670 15450 8676
rect 15326 8636 15338 8670
rect 15438 8636 15450 8670
rect 15326 8630 15450 8636
rect 15506 8598 15561 8750
rect 15726 8670 15850 8676
rect 15726 8636 15738 8670
rect 15838 8636 15850 8670
rect 15726 8630 15850 8636
rect 15906 8598 15961 8750
rect 16815 8792 16890 8872
rect 17189 8792 17270 8879
rect 16815 8749 17270 8792
rect 16126 8670 16250 8676
rect 16126 8636 16138 8670
rect 16238 8636 16250 8670
rect 16126 8630 16250 8636
rect 16526 8670 16650 8676
rect 16526 8636 16538 8670
rect 16638 8636 16650 8670
rect 16526 8630 16650 8636
rect 16815 8598 16870 8749
rect 16926 8670 17050 8676
rect 16926 8636 16938 8670
rect 17038 8636 17050 8670
rect 16926 8630 17050 8636
rect 17215 8598 17270 8749
rect 17326 8670 17450 8676
rect 17326 8636 17338 8670
rect 17438 8636 17450 8670
rect 17326 8630 17450 8636
rect 17615 8598 17670 8990
rect 17726 8670 17850 8676
rect 17726 8636 17738 8670
rect 17838 8636 17850 8670
rect 17726 8630 17850 8636
rect 18126 8670 18250 8676
rect 18126 8636 18138 8670
rect 18238 8636 18250 8670
rect 18126 8630 18250 8636
rect 14470 8586 14516 8598
rect 14470 7590 14476 8586
rect 14510 7590 14516 8586
rect 14470 7578 14516 7590
rect 14660 8586 14706 8598
rect 14660 7590 14666 8586
rect 14700 7590 14706 8586
rect 14660 7578 14706 7590
rect 14870 8586 14916 8598
rect 14870 7590 14876 8586
rect 14910 7590 14916 8586
rect 14870 7578 14916 7590
rect 15060 8586 15161 8598
rect 15060 7590 15066 8586
rect 15100 7590 15161 8586
rect 15060 7578 15161 7590
rect 15270 8586 15316 8598
rect 15270 7590 15276 8586
rect 15310 7590 15316 8586
rect 15270 7578 15316 7590
rect 15460 8586 15561 8598
rect 15460 7590 15466 8586
rect 15500 7590 15561 8586
rect 15460 7578 15561 7590
rect 15670 8586 15716 8598
rect 15670 7590 15676 8586
rect 15710 7590 15716 8586
rect 15670 7578 15716 7590
rect 15860 8586 15961 8598
rect 15860 7590 15866 8586
rect 15900 7590 15961 8586
rect 15860 7578 15961 7590
rect 16070 8586 16116 8598
rect 16070 7590 16076 8586
rect 16110 7590 16116 8586
rect 16070 7578 16116 7590
rect 16260 8586 16516 8598
rect 16260 7590 16266 8586
rect 16300 7590 16476 8586
rect 16510 7590 16516 8586
rect 16260 7578 16516 7590
rect 16660 8586 16706 8598
rect 16660 7590 16666 8586
rect 16700 7590 16706 8586
rect 16660 7578 16706 7590
rect 16815 8586 16916 8598
rect 16815 7590 16876 8586
rect 16910 7590 16916 8586
rect 16815 7578 16916 7590
rect 17060 8586 17106 8598
rect 17060 7590 17066 8586
rect 17100 7590 17106 8586
rect 17060 7578 17106 7590
rect 17215 8586 17316 8598
rect 17215 7590 17276 8586
rect 17310 7590 17316 8586
rect 17215 7578 17316 7590
rect 17460 8586 17506 8598
rect 17460 7590 17466 8586
rect 17500 7590 17506 8586
rect 17460 7578 17506 7590
rect 17615 8586 17716 8598
rect 17615 7590 17676 8586
rect 17710 7590 17716 8586
rect 17615 7578 17716 7590
rect 17860 8586 17906 8598
rect 17860 7590 17866 8586
rect 17900 7590 17906 8586
rect 17860 7578 17906 7590
rect 18070 8586 18116 8598
rect 18070 7590 18076 8586
rect 18110 7590 18116 8586
rect 18070 7578 18116 7590
rect 18260 8586 18306 8598
rect 18260 7590 18266 8586
rect 18300 7590 18306 8586
rect 18260 7578 18306 7590
rect 14526 7540 14650 7546
rect 14526 7506 14538 7540
rect 14638 7506 14650 7540
rect 14526 7500 14650 7506
rect 14926 7540 15050 7546
rect 14926 7506 14938 7540
rect 15038 7512 15050 7540
rect 15326 7540 15450 7546
rect 15326 7512 15338 7540
rect 15038 7506 15338 7512
rect 15438 7512 15450 7540
rect 15726 7540 15850 7546
rect 15726 7512 15738 7540
rect 15438 7506 15738 7512
rect 15838 7512 15850 7540
rect 16126 7540 16250 7546
rect 16126 7512 16138 7540
rect 15838 7506 16138 7512
rect 16238 7512 16250 7540
rect 16356 7512 16415 7578
rect 16526 7540 16650 7546
rect 16526 7512 16538 7540
rect 16238 7506 16538 7512
rect 16638 7512 16650 7540
rect 16926 7540 17050 7546
rect 16926 7512 16938 7540
rect 16638 7506 16938 7512
rect 17038 7512 17050 7540
rect 17326 7540 17450 7546
rect 17326 7512 17338 7540
rect 17038 7506 17338 7512
rect 17438 7512 17450 7540
rect 17726 7540 17850 7546
rect 17726 7512 17738 7540
rect 17438 7506 17738 7512
rect 17838 7506 17850 7540
rect 14926 7442 17850 7506
rect 18126 7540 18250 7546
rect 18126 7506 18138 7540
rect 18238 7506 18250 7540
rect 18126 7500 18250 7506
rect 16316 7327 16465 7442
rect 16311 7296 16465 7327
rect 16311 7117 18938 7296
rect -726 5482 18815 6140
<< via1 >>
rect 1151 18558 1234 18718
rect 548 17358 649 17606
rect -320 15349 -55 15546
rect 1148 16191 1231 16351
rect 2954 16051 3006 17963
rect 11162 17720 12344 17945
rect 9084 16473 9786 16574
rect 9084 16379 9594 16473
rect 9594 16379 9786 16473
rect 3598 15391 3653 15673
rect 16114 17288 16166 17434
rect 17510 17288 17562 17434
rect 17590 17078 17646 17276
rect 16114 16918 16166 17064
rect 17510 16918 17562 17064
rect 15770 16308 15970 16370
rect 17234 16438 17336 16562
rect 749 14940 826 14996
rect 1894 14940 1971 14996
rect 9274 15242 9372 15246
rect 9274 15194 9371 15242
rect 9371 15194 9372 15242
rect 9645 15242 9743 15246
rect 9645 15194 9646 15242
rect 9646 15194 9743 15242
rect 2698 14566 2788 14786
rect 2055 13102 2220 13608
rect 2699 12164 2789 12384
rect 9291 14761 9354 14829
rect 9663 14761 9726 14829
rect 9274 13576 9372 13580
rect 9274 13528 9371 13576
rect 9371 13528 9372 13576
rect 9645 13576 9743 13580
rect 9645 13528 9646 13576
rect 9646 13528 9743 13576
rect 9291 13095 9354 13163
rect 9663 13095 9726 13163
rect 3598 11300 3653 11582
rect 2420 8504 2762 9116
rect 2954 8995 3006 10907
rect 9274 11910 9372 11914
rect 9274 11862 9371 11910
rect 9371 11862 9372 11910
rect 9645 11910 9743 11914
rect 9645 11862 9646 11910
rect 9646 11862 9743 11910
rect 9291 11429 9354 11497
rect 9663 11429 9726 11497
rect 9274 10244 9372 10248
rect 9274 10196 9371 10244
rect 9371 10196 9372 10244
rect 9645 10244 9743 10248
rect 9645 10196 9646 10244
rect 9646 10196 9743 10244
rect 3874 8735 4110 8827
rect -291 7595 59 7832
rect 4854 7246 5270 9676
rect 9291 9763 9354 9831
rect 9663 9763 9726 9831
rect 9274 8578 9372 8582
rect 9274 8530 9371 8578
rect 9371 8530 9372 8578
rect 9645 8578 9743 8582
rect 9645 8530 9646 8578
rect 9646 8530 9743 8578
rect 9291 8097 9354 8165
rect 9663 8097 9726 8165
rect 16258 12664 16384 12815
rect 14975 12442 15349 12532
rect 14431 12043 14693 12225
rect 14872 10673 14880 11536
rect 14880 10673 14924 11536
rect 15078 11092 15159 11768
rect 14867 9519 14880 10382
rect 14880 9519 14919 10382
rect 16562 12264 16633 12382
rect 16750 11266 16829 11549
rect 17124 10640 17596 10942
rect 17058 9153 17230 9283
rect 15580 8792 15879 8879
rect 16890 8792 17189 8879
<< metal2 >>
rect 1137 18718 1251 18753
rect 1137 18558 1151 18718
rect 1234 18558 1251 18718
rect 1137 18527 1251 18558
rect 530 17606 680 17674
rect 530 17358 548 17606
rect 649 17358 680 17606
rect 530 17298 680 17358
rect 594 16865 671 17298
rect 872 16865 982 16867
rect 594 16771 982 16865
rect -345 15546 -23 15580
rect -345 15542 -320 15546
rect -346 15349 -320 15542
rect -55 15349 -23 15546
rect -346 15320 -23 15349
rect -346 7893 -202 15320
rect 872 15240 982 16771
rect 1155 16384 1230 18527
rect 2934 17963 3024 18046
rect 12233 17992 12413 20748
rect 1135 16351 1249 16384
rect 1135 16191 1148 16351
rect 1231 16191 1249 16351
rect 1135 16158 1249 16191
rect 2934 16051 2954 17963
rect 3006 16051 3024 17963
rect 11103 17945 12417 17992
rect 11103 17720 11162 17945
rect 12344 17720 12417 17945
rect 11103 17676 12417 17720
rect 16104 17434 16206 17446
rect 16104 17288 16114 17434
rect 16166 17288 16206 17434
rect 16104 17276 16206 17288
rect 17470 17434 17660 17446
rect 17470 17288 17510 17434
rect 17562 17288 17660 17434
rect 17470 17276 17660 17288
rect 16104 17076 16160 17276
rect 17516 17078 17590 17276
rect 17646 17078 17660 17276
rect 17516 17076 17660 17078
rect 16104 17064 16206 17076
rect 16104 16918 16114 17064
rect 16166 16918 16206 17064
rect 16104 16906 16206 16918
rect 17470 17064 17660 17076
rect 17470 16918 17510 17064
rect 17562 16918 17660 17064
rect 17470 16906 17660 16918
rect 9010 16574 9850 16628
rect 9010 16379 9084 16574
rect 9786 16379 9850 16574
rect 17210 16562 17362 16584
rect 17210 16438 17234 16562
rect 17336 16438 17362 16562
rect 17210 16420 17362 16438
rect 9010 16343 9850 16379
rect 15770 16370 16058 16396
rect 871 15138 2809 15240
rect 711 14996 864 15020
rect 711 14940 749 14996
rect 826 14989 864 14996
rect 1856 15001 2009 15020
rect 1856 14996 2534 15001
rect 1856 14989 1894 14996
rect 826 14942 1894 14989
rect 826 14940 864 14942
rect 711 14923 864 14940
rect 1856 14940 1894 14942
rect 1971 14940 2534 14996
rect 1856 14925 2534 14940
rect 1856 14923 2009 14925
rect 1854 13611 2285 13685
rect 1854 13072 1893 13611
rect 2228 13072 2285 13611
rect 1854 13005 2285 13072
rect 2420 10888 2534 14925
rect 2679 14786 2809 15138
rect 2679 14566 2698 14786
rect 2788 14566 2809 14786
rect 2679 12446 2809 14566
rect 2679 12384 2810 12446
rect 2679 12246 2699 12384
rect 2680 12164 2699 12246
rect 2789 12164 2810 12384
rect 2680 12104 2810 12164
rect 2934 10907 3024 16051
rect 9052 15789 9178 16343
rect 15970 16308 16058 16370
rect 15770 16278 16058 16308
rect 16000 16184 16058 16278
rect 17260 16184 17362 16420
rect 16000 16114 17362 16184
rect 16482 15937 16626 16114
rect 16482 15844 18576 15937
rect 8713 15746 9178 15789
rect 8712 15732 9178 15746
rect 3593 15673 3658 15681
rect 3593 15391 3598 15673
rect 3653 15391 3658 15673
rect 3593 11582 3658 15391
rect 8712 15284 8852 15732
rect 16483 15706 18576 15844
rect 8712 15264 9402 15284
rect 8712 15250 9436 15264
rect 8712 15194 9274 15250
rect 9377 15194 9436 15250
rect 8712 15179 9436 15194
rect 9581 15263 10287 15264
rect 9581 15250 10308 15263
rect 9581 15194 9640 15250
rect 9743 15194 10308 15250
rect 9581 15179 10308 15194
rect 8712 15170 9402 15179
rect 9271 14837 9376 14851
rect 9641 14837 9746 14851
rect 9271 14829 9746 14837
rect 9271 14761 9291 14829
rect 9354 14761 9663 14829
rect 9726 14761 9746 14829
rect 9271 14759 9746 14761
rect 9271 14744 9376 14759
rect 9641 14744 9746 14759
rect 9249 13584 9436 13598
rect 9249 13528 9274 13584
rect 9377 13528 9436 13584
rect 9249 13513 9436 13528
rect 9581 13584 9768 13598
rect 9581 13528 9640 13584
rect 9743 13528 9768 13584
rect 9581 13513 9768 13528
rect 9271 13172 9376 13185
rect 8711 13163 9376 13172
rect 8711 13095 9291 13163
rect 9354 13095 9376 13163
rect 8711 13087 9376 13095
rect 8711 11932 8823 13087
rect 9271 13078 9376 13087
rect 9641 13180 9746 13185
rect 10204 13180 10308 15179
rect 9641 13163 10308 13180
rect 9641 13095 9663 13163
rect 9726 13095 10308 13163
rect 9641 13078 9746 13095
rect 16218 12815 16424 12869
rect 16218 12664 16258 12815
rect 16384 12664 16424 12815
rect 16218 12626 16424 12664
rect 14899 12554 15418 12555
rect 16252 12554 16395 12626
rect 14899 12532 16395 12554
rect 14899 12442 14975 12532
rect 15349 12442 16395 12532
rect 14899 12423 16395 12442
rect 14899 12422 16331 12423
rect 16532 12382 16664 12421
rect 16532 12300 16562 12382
rect 14732 12298 16562 12300
rect 14340 12264 16562 12298
rect 16633 12300 16664 12382
rect 16633 12264 16822 12300
rect 14340 12241 16822 12264
rect 14340 12226 14965 12241
rect 14340 12225 14787 12226
rect 14340 12043 14431 12225
rect 14693 12043 14787 12225
rect 14340 11971 14787 12043
rect 14911 12044 14965 12226
rect 15171 12226 16822 12241
rect 15171 12044 15228 12226
rect 14911 11997 15228 12044
rect 8711 11918 9436 11932
rect 8711 11862 9274 11918
rect 9377 11862 9436 11918
rect 8711 11847 9436 11862
rect 9581 11931 10287 11932
rect 9581 11918 10308 11931
rect 9581 11862 9640 11918
rect 9743 11862 10308 11918
rect 9581 11847 10308 11862
rect 3593 11300 3598 11582
rect 3653 11300 3658 11582
rect 9271 11497 9376 11519
rect 9271 11429 9291 11497
rect 9354 11429 9376 11497
rect 9271 11412 9376 11429
rect 9641 11497 9746 11519
rect 9641 11429 9663 11497
rect 9726 11429 9746 11497
rect 9641 11412 9746 11429
rect 3593 11292 3658 11300
rect 2420 10887 2703 10888
rect 2934 10887 2954 10907
rect 2420 10674 2954 10887
rect 2442 10673 2954 10674
rect 2639 10577 2954 10673
rect 2376 9116 2814 9166
rect 2376 8504 2420 9116
rect 2762 8504 2814 9116
rect 2934 8995 2954 10577
rect 3006 8995 3024 10907
rect 9249 10252 9436 10266
rect 9249 10196 9274 10252
rect 9377 10196 9436 10252
rect 9249 10181 9436 10196
rect 9581 10252 9768 10266
rect 9581 10196 9640 10252
rect 9743 10196 9768 10252
rect 9581 10181 9768 10196
rect 9271 9844 9376 9853
rect 8711 9831 9376 9844
rect 8711 9763 9291 9831
rect 9354 9763 9376 9831
rect 2934 8832 3024 8995
rect 4766 9676 5354 9760
rect 3786 8832 4178 8881
rect 2934 8827 4178 8832
rect 2934 8737 3874 8827
rect 3786 8735 3874 8737
rect 4110 8735 4178 8827
rect 3786 8679 4178 8735
rect 2376 8454 2814 8504
rect -347 7832 116 7893
rect -347 7595 -291 7832
rect 59 7595 116 7832
rect -347 7545 116 7595
rect 2502 7782 2712 8454
rect 2502 7781 2864 7782
rect 4766 7781 4854 9676
rect 2502 7246 4854 7781
rect 5270 7246 5354 9676
rect 8711 9759 9376 9763
rect 8711 8600 8823 9759
rect 9271 9746 9376 9759
rect 9641 9848 9746 9853
rect 10204 9848 10308 11847
rect 15043 11768 15198 11814
rect 14840 11536 14952 11566
rect 14840 10673 14872 11536
rect 14924 10696 14952 11536
rect 15043 11092 15078 11768
rect 15159 11758 15198 11768
rect 15159 11696 15335 11758
rect 15285 11098 15335 11696
rect 16722 11583 16822 12226
rect 16722 11549 16857 11583
rect 16722 11266 16750 11549
rect 16829 11266 16857 11549
rect 16722 11238 16857 11266
rect 15159 11092 15335 11098
rect 15043 11050 15335 11092
rect 17058 10942 17654 10988
rect 14924 10673 15170 10696
rect 14840 10636 15170 10673
rect 14902 10418 15170 10636
rect 17058 10640 17124 10942
rect 17596 10640 17654 10942
rect 17058 10592 17654 10640
rect 9641 9831 10308 9848
rect 9641 9763 9663 9831
rect 9726 9763 10308 9831
rect 14840 10382 15170 10418
rect 9641 9746 9746 9763
rect 14840 9519 14867 10382
rect 14919 10339 15170 10382
rect 14919 9519 14952 10339
rect 14840 9488 14952 9519
rect 15035 8921 15170 10339
rect 17027 9283 17270 9317
rect 17027 9153 17058 9283
rect 17230 9153 17270 9283
rect 15035 8920 15633 8921
rect 17027 8920 17270 9153
rect 15035 8900 15961 8920
rect 15036 8879 15961 8900
rect 15036 8837 15580 8879
rect 15506 8792 15580 8837
rect 15879 8792 15961 8879
rect 15506 8750 15961 8792
rect 16815 8879 17270 8920
rect 16815 8792 16890 8879
rect 17189 8792 17270 8879
rect 16815 8749 17270 8792
rect 8711 8586 9436 8600
rect 8711 8530 9274 8586
rect 9377 8530 9436 8586
rect 8711 8515 9436 8530
rect 9581 8586 10289 8600
rect 9581 8530 9640 8586
rect 9743 8530 10289 8586
rect 9581 8515 10289 8530
rect 9271 8178 9376 8187
rect 9271 8165 9542 8178
rect 9271 8097 9291 8165
rect 9354 8126 9542 8165
rect 9354 8097 9376 8126
rect 9271 8080 9376 8097
rect 9462 7384 9542 8126
rect 9641 8165 9746 8187
rect 9641 8097 9663 8165
rect 9726 8097 9746 8165
rect 9641 8080 9746 8097
rect 10198 7384 10289 8515
rect 9462 7320 10289 7384
rect 2502 7243 5354 7246
rect 2502 7242 2842 7243
rect 4766 7166 5354 7243
<< via2 >>
rect 1893 13608 2228 13611
rect 1893 13102 2055 13608
rect 2055 13102 2220 13608
rect 2220 13102 2228 13608
rect 1893 13072 2228 13102
rect 9274 15246 9377 15250
rect 9274 15194 9372 15246
rect 9372 15194 9377 15246
rect 9640 15246 9743 15250
rect 9640 15194 9645 15246
rect 9645 15194 9743 15246
rect 9291 14761 9354 14829
rect 9663 14761 9726 14829
rect 9274 13580 9377 13584
rect 9274 13528 9372 13580
rect 9372 13528 9377 13580
rect 9640 13580 9743 13584
rect 9640 13528 9645 13580
rect 9645 13528 9743 13580
rect 9291 13095 9354 13163
rect 9663 13095 9726 13163
rect 14965 12044 15171 12241
rect 9274 11914 9377 11918
rect 9274 11862 9372 11914
rect 9372 11862 9377 11914
rect 9640 11914 9743 11918
rect 9640 11862 9645 11914
rect 9645 11862 9743 11914
rect 9291 11429 9354 11497
rect 9663 11429 9726 11497
rect 9274 10248 9377 10252
rect 9274 10196 9372 10248
rect 9372 10196 9377 10248
rect 9640 10248 9743 10252
rect 9640 10196 9645 10248
rect 9645 10196 9743 10248
rect 9291 9763 9354 9831
rect 15088 11098 15159 11696
rect 15159 11098 15285 11696
rect 17124 10640 17596 10942
rect 9663 9763 9726 9831
rect 9274 8582 9377 8586
rect 9274 8530 9372 8582
rect 9372 8530 9377 8582
rect 9640 8582 9743 8586
rect 9640 8530 9645 8582
rect 9645 8530 9743 8582
rect 9291 8097 9354 8165
rect 9663 8097 9726 8165
<< metal3 >>
rect 9249 15250 9436 15264
rect 9249 15194 9274 15250
rect 9377 15194 9436 15250
rect 9249 15179 9436 15194
rect 9581 15250 9768 15264
rect 9581 15194 9640 15250
rect 9743 15194 9768 15250
rect 9581 15179 9768 15194
rect 9247 14841 9400 14877
rect 8709 14829 9400 14841
rect 8709 14761 9291 14829
rect 9354 14761 9400 14829
rect 8709 14756 9400 14761
rect 1854 13611 2285 13685
rect 1854 13301 1893 13611
rect -475 13072 1893 13301
rect 2228 13072 2285 13611
rect 8709 13599 8821 14756
rect 9247 14726 9400 14756
rect 9617 14829 9770 14877
rect 9617 14761 9663 14829
rect 9726 14761 9770 14829
rect 9617 14726 9770 14761
rect 8709 13598 9397 13599
rect 8709 13584 9436 13598
rect 8709 13528 9274 13584
rect 9377 13528 9436 13584
rect 8709 13514 9436 13528
rect 9249 13513 9436 13514
rect 9581 13597 10287 13598
rect 9581 13584 10308 13597
rect 9581 13528 9640 13584
rect 9743 13528 10308 13584
rect 9581 13513 10308 13528
rect -475 13014 2285 13072
rect 9247 13163 9400 13211
rect 9247 13095 9291 13163
rect 9354 13095 9400 13163
rect 9247 13060 9400 13095
rect 9617 13163 9770 13211
rect 9617 13095 9663 13163
rect 9726 13095 9770 13163
rect 9617 13060 9770 13095
rect -475 10504 -281 13014
rect 1854 13005 2285 13014
rect 9249 11918 9436 11932
rect 9249 11862 9274 11918
rect 9377 11862 9436 11918
rect 9249 11847 9436 11862
rect 9581 11918 9768 11932
rect 9581 11862 9640 11918
rect 9743 11862 9768 11918
rect 9581 11847 9768 11862
rect 9247 11504 9400 11545
rect 8708 11497 9400 11504
rect 8708 11429 9291 11497
rect 9354 11429 9400 11497
rect 8708 11419 9400 11429
rect -475 10226 64 10504
rect -120 9515 64 10226
rect 8708 10266 8820 11419
rect 9247 11394 9400 11419
rect 9617 11514 9770 11545
rect 10204 11514 10308 13513
rect 14911 12241 15228 12300
rect 14911 12044 14965 12241
rect 15171 12044 15228 12241
rect 14911 11997 15228 12044
rect 15496 12177 16668 12205
rect 9617 11497 10308 11514
rect 9617 11429 9663 11497
rect 9726 11429 10308 11497
rect 15043 11696 15335 11758
rect 9617 11394 9770 11429
rect 15043 11098 15088 11696
rect 15285 11098 15335 11696
rect 15043 11050 15335 11098
rect 8708 10252 9436 10266
rect 8708 10196 9274 10252
rect 9377 10196 9436 10252
rect 8708 10181 9436 10196
rect 9581 10265 10287 10266
rect 9581 10252 10308 10265
rect 9581 10196 9640 10252
rect 9743 10196 10308 10252
rect 9581 10181 10308 10196
rect 9247 9831 9400 9879
rect 9247 9763 9291 9831
rect 9354 9763 9400 9831
rect 9247 9728 9400 9763
rect 9617 9831 9770 9879
rect 9617 9763 9663 9831
rect 9726 9763 9770 9831
rect 9617 9728 9770 9763
rect -120 9174 769 9515
rect -1074 8423 769 9174
rect 9249 8586 9436 8600
rect 9249 8530 9274 8586
rect 9377 8530 9436 8586
rect 9249 8515 9436 8530
rect 9581 8586 9768 8600
rect 9581 8530 9640 8586
rect 9743 8530 9768 8586
rect 9581 8515 9768 8530
rect -120 8087 769 8423
rect 9247 8165 9400 8213
rect 9247 8097 9291 8165
rect 9354 8097 9400 8165
rect 9247 8062 9400 8097
rect 9617 8182 9770 8213
rect 10204 8182 10308 10181
rect 15210 9016 15335 11050
rect 15496 9153 16584 12177
rect 16648 9153 16668 12177
rect 17058 10942 17654 10988
rect 17058 10640 17124 10942
rect 17596 10640 17654 10942
rect 17058 10592 17654 10640
rect 15496 9125 16668 9153
rect 18158 9016 18870 9125
rect 15210 8894 18870 9016
rect 15210 8886 18243 8894
rect 9617 8165 10308 8182
rect 9617 8097 9663 8165
rect 9726 8097 10308 8165
rect 9617 8062 9770 8097
<< via3 >>
rect 14965 12044 15171 12241
rect 16584 9153 16648 12177
rect 17124 10640 17596 10942
<< mimcap >>
rect 15536 12125 16336 12165
rect 15536 9205 15576 12125
rect 16296 9205 16336 12125
rect 15536 9165 16336 9205
<< mimcapcontact >>
rect 15576 9205 16296 12125
<< metal4 >>
rect 14911 12241 15228 12300
rect 14911 12044 14965 12241
rect 15171 12126 15228 12241
rect 16568 12177 16664 12193
rect 15171 12125 16297 12126
rect 15171 12044 15576 12125
rect 14911 11997 15576 12044
rect 15575 9205 15576 11997
rect 16296 9205 16297 12125
rect 15575 9204 16297 9205
rect 16568 9153 16584 12177
rect 16648 10914 16664 12177
rect 17058 10942 17654 10988
rect 17058 10914 17124 10942
rect 16648 10654 17124 10914
rect 16648 9153 16664 10654
rect 17058 10640 17124 10654
rect 17596 10640 17654 10942
rect 17058 10592 17654 10640
rect 16568 9137 16664 9153
<< labels >>
flabel metal2 12262 20580 12382 20694 0 FreeSans 3200 90 0 0 ring_out
port 0 nsew
flabel metal1 13290 20582 13410 20696 0 FreeSans 3200 90 0 0 dd_02
port 1 nsew
flabel metal2 17886 15766 18006 15880 0 FreeSans 3200 0 0 0 vref
port 2 nsew
flabel metal1 18374 10724 18494 10838 0 FreeSans 3200 0 0 0 ldo_out
port 3 nsew
flabel metal1 18674 10062 18748 10150 0 FreeSans 3200 0 0 0 ldo_vs
port 4 nsew
flabel metal3 18678 8958 18752 9046 0 FreeSans 3200 0 0 0 ldo_vb
port 5 nsew
flabel metal1 18716 7170 18790 7258 0 FreeSans 3200 0 0 0 ldo_iref
port 6 nsew
flabel metal1 18374 5776 18448 5864 0 FreeSans 3200 0 0 0 dd_01
port 7 nsew
flabel locali -718 6724 -526 6906 0 FreeSans 3200 0 0 0 ss
port 8 nsew
flabel metal3 -840 8674 -648 8856 0 FreeSans 3200 0 0 0 iref
port 9 nsew
flabel metal2 16020 16122 16088 16170 0 FreeSans 1600 0 0 0 vref01_0.VREF
flabel metal1 15956 17472 16024 17520 0 FreeSans 1600 0 0 0 vref01_0.DD
flabel locali 17734 16464 17802 16512 0 FreeSans 1600 0 0 0 vref01_0.SS
flabel locali 6256 15787 6604 16039 0 FreeSans 1600 0 0 0 ring_100mV_0.SS
flabel metal1 11058 15897 11264 16087 0 FreeSans 1600 0 0 0 ring_100mV_0.DD
flabel space 11690 17761 11896 17951 0 FreeSans 1600 0 0 0 ring_100mV_0.OUT
flabel metal1 11994 17800 12122 17904 0 FreeSans 1600 0 0 0 ring_100mV_0.ring_100mV_buffer_0.OUT
flabel metal2 9695 16490 9823 16594 0 FreeSans 1600 0 0 0 ring_100mV_0.ring_100mV_buffer_0.IN
flabel viali 10600 16465 10728 16569 0 FreeSans 1600 0 0 0 ring_100mV_0.ring_100mV_buffer_0.DD
flabel locali 5482 16153 5610 16257 0 FreeSans 1600 0 0 0 ring_100mV_0.ring_100mV_buffer_0.SS
rlabel metal1 10239 9318 10314 9382 7 ring_100mV_0.mdls_inv_9.IN
rlabel locali 11191 10647 11266 10711 7 ring_100mV_0.mdls_inv_9.SS
rlabel locali 9614 10593 9652 10627 7 ring_100mV_0.mdls_inv_9.DD
rlabel metal1 11785 10553 11829 10592 7 ring_100mV_0.mdls_inv_9.OUT
rlabel metal1 8703 9318 8778 9382 3 ring_100mV_0.mdls_inv_8.IN
rlabel locali 7751 10647 7826 10711 3 ring_100mV_0.mdls_inv_8.SS
rlabel locali 9365 10593 9403 10627 3 ring_100mV_0.mdls_inv_8.DD
rlabel metal1 7188 10553 7232 10592 3 ring_100mV_0.mdls_inv_8.OUT
rlabel metal1 10239 10984 10314 11048 7 ring_100mV_0.mdls_inv_7.IN
rlabel locali 11191 12313 11266 12377 7 ring_100mV_0.mdls_inv_7.SS
rlabel locali 9614 12259 9652 12293 7 ring_100mV_0.mdls_inv_7.DD
rlabel metal1 11785 12219 11829 12258 7 ring_100mV_0.mdls_inv_7.OUT
rlabel metal1 8703 10984 8778 11048 3 ring_100mV_0.mdls_inv_6.IN
rlabel locali 7751 12313 7826 12377 3 ring_100mV_0.mdls_inv_6.SS
rlabel locali 9365 12259 9403 12293 3 ring_100mV_0.mdls_inv_6.DD
rlabel metal1 7188 12219 7232 12258 3 ring_100mV_0.mdls_inv_6.OUT
rlabel metal1 10239 12650 10314 12714 7 ring_100mV_0.mdls_inv_5.IN
rlabel locali 11191 13979 11266 14043 7 ring_100mV_0.mdls_inv_5.SS
rlabel locali 9614 13925 9652 13959 7 ring_100mV_0.mdls_inv_5.DD
rlabel metal1 11785 13885 11829 13924 7 ring_100mV_0.mdls_inv_5.OUT
rlabel metal1 8703 12650 8778 12714 3 ring_100mV_0.mdls_inv_4.IN
rlabel locali 7751 13979 7826 14043 3 ring_100mV_0.mdls_inv_4.SS
rlabel locali 9365 13925 9403 13959 3 ring_100mV_0.mdls_inv_4.DD
rlabel metal1 7188 13885 7232 13924 3 ring_100mV_0.mdls_inv_4.OUT
rlabel metal1 8703 14316 8778 14380 3 ring_100mV_0.mdls_inv_3.IN
rlabel locali 7751 15645 7826 15709 3 ring_100mV_0.mdls_inv_3.SS
rlabel locali 9365 15591 9403 15625 3 ring_100mV_0.mdls_inv_3.DD
rlabel metal1 7188 15551 7232 15590 3 ring_100mV_0.mdls_inv_3.OUT
rlabel metal1 10239 14316 10314 14380 7 ring_100mV_0.mdls_inv_2.IN
rlabel locali 11191 15645 11266 15709 7 ring_100mV_0.mdls_inv_2.SS
rlabel locali 9614 15591 9652 15625 7 ring_100mV_0.mdls_inv_2.DD
rlabel metal1 11785 15551 11829 15590 7 ring_100mV_0.mdls_inv_2.OUT
rlabel metal1 8703 7652 8778 7716 3 ring_100mV_0.mdls_inv_1.IN
rlabel locali 7751 8981 7826 9045 3 ring_100mV_0.mdls_inv_1.SS
rlabel locali 9365 8927 9403 8961 3 ring_100mV_0.mdls_inv_1.DD
rlabel metal1 7188 8887 7232 8926 3 ring_100mV_0.mdls_inv_1.OUT
rlabel metal1 10239 7652 10314 7716 7 ring_100mV_0.mdls_inv_0.IN
rlabel locali 11191 8981 11266 9045 7 ring_100mV_0.mdls_inv_0.SS
rlabel locali 9614 8927 9652 8961 7 ring_100mV_0.mdls_inv_0.DD
rlabel metal1 11785 8887 11829 8926 7 ring_100mV_0.mdls_inv_0.OUT
flabel metal1 16352 7712 16428 7800 0 FreeSans 1600 0 0 0 ldo_0.Iref
flabel locali 14614 8942 14690 9030 0 FreeSans 1600 0 0 0 ldo_0.SS
flabel metal3 18264 8932 18438 9064 0 FreeSans 1600 0 0 0 ldo_0.VB
flabel metal1 18490 10082 18540 10136 0 FreeSans 1600 0 0 0 ldo_0.VS
flabel metal1 18084 10672 18284 10848 0 FreeSans 1600 0 0 0 ldo_0.OUT
flabel metal1 18376 13500 18468 13616 0 FreeSans 1600 0 0 0 ldo_0.DD
flabel metal2 3910 7478 4140 7682 0 FreeSans 1600 0 0 0 iref_2nA_0.DD
flabel metal3 210 8766 440 8970 0 FreeSans 1600 0 0 0 iref_2nA_0.IREF
flabel locali 570 19250 718 19414 0 FreeSans 1600 0 0 0 iref_2nA_0.SS
flabel locali 2155 9785 2233 9863 0 FreeSans 1600 0 0 0 iref_2nA_0.iref_2nA_vref_0.DD
flabel locali 2477 11747 2551 11833 0 FreeSans 1600 0 0 0 iref_2nA_0.iref_2nA_vref_0.SS
flabel metal1 69 11759 143 11845 0 FreeSans 1600 0 0 0 iref_2nA_0.iref_2nA_vref_0.VREF
rlabel metal2 2680 10636 2815 10846 5 iref_2nA_0.iref_2nA_mirrors_0.Ip2
rlabel metal1 2610 13444 2660 13517 5 iref_2nA_0.iref_2nA_mirrors_0.Iref
rlabel metal1 842 17371 892 17444 5 iref_2nA_0.iref_2nA_mirrors_0.Vg
rlabel metal2 1156 18591 1206 18664 5 iref_2nA_0.iref_2nA_mirrors_0.Ip1
rlabel locali 112 19274 238 19379 5 iref_2nA_0.iref_2nA_mirrors_0.SS
rlabel locali 2579 8468 2667 8542 5 iref_2nA_0.iref_2nA_mirrors_0.DD
rlabel metal1 -302 14877 -260 14935 7 iref_2nA_0.iref_2nA_igenerator_0.Vg
rlabel metal1 1132 14685 1174 14743 7 iref_2nA_0.iref_2nA_igenerator_0.Ip1
rlabel metal1 718 14685 760 14743 7 iref_2nA_0.iref_2nA_igenerator_0.Ip2
rlabel locali 550 13599 592 13657 7 iref_2nA_0.iref_2nA_igenerator_0.SS
rlabel metal1 346 13579 388 13637 7 iref_2nA_0.iref_2nA_igenerator_0.VCTAT
<< end >>

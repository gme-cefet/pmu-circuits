magic
tech sky130A
magscale 1 2
timestamp 1695321174
<< error_p >>
rect 6234 7884 6249 7912
rect 6262 7690 6277 7884
<< error_s >>
rect 8071 8180 9345 8230
rect 9507 8180 10799 8230
rect 8358 8168 8359 8179
rect 8670 8168 8671 8179
rect 8982 8168 8983 8179
rect 9294 8168 9295 8179
rect 9812 8168 9813 8179
rect 10124 8168 10125 8179
rect 10436 8168 10437 8179
rect 10748 8168 10749 8179
rect 8202 8126 8203 8137
rect 8369 8134 8370 8168
rect 8514 8126 8515 8137
rect 8681 8134 8682 8168
rect 8826 8126 8827 8137
rect 8993 8134 8994 8168
rect 9138 8126 9139 8137
rect 9305 8134 9306 8168
rect 9656 8126 9657 8137
rect 9823 8134 9824 8168
rect 9968 8126 9969 8137
rect 10135 8134 10136 8168
rect 10280 8126 10281 8137
rect 10447 8134 10448 8168
rect 10592 8126 10593 8137
rect 10759 8134 10760 8168
rect 8213 8092 8214 8126
rect 8358 8100 8359 8111
rect 8202 8058 8203 8069
rect 8369 8066 8370 8100
rect 8525 8092 8526 8126
rect 8670 8100 8671 8111
rect 8514 8058 8515 8069
rect 8681 8066 8682 8100
rect 8837 8092 8838 8126
rect 8982 8100 8983 8111
rect 8826 8058 8827 8069
rect 8993 8066 8994 8100
rect 9149 8092 9150 8126
rect 9294 8100 9295 8111
rect 9138 8058 9139 8069
rect 8213 8024 8214 8058
rect 8358 8032 8359 8043
rect 8202 7990 8203 8001
rect 8369 7998 8370 8032
rect 8525 8024 8526 8058
rect 8670 8032 8671 8043
rect 8514 7990 8515 8001
rect 8681 7998 8682 8032
rect 8837 8024 8838 8058
rect 8982 8032 8983 8043
rect 8826 7990 8827 8001
rect 8993 7998 8994 8032
rect 9149 8024 9150 8058
rect 9138 7990 9139 8001
rect 8213 7956 8214 7990
rect 8358 7964 8359 7975
rect 8202 7922 8203 7933
rect 8369 7930 8370 7964
rect 8525 7956 8526 7990
rect 8670 7964 8671 7975
rect 8514 7922 8515 7933
rect 8681 7930 8682 7964
rect 8837 7956 8838 7990
rect 8982 7964 8983 7975
rect 8826 7922 8827 7933
rect 8993 7930 8994 7964
rect 9149 7956 9150 7990
rect 9138 7922 9139 7933
rect 8213 7888 8214 7922
rect 8525 7888 8526 7922
rect 8837 7888 8838 7922
rect 9149 7888 9150 7922
rect 9269 7880 9270 8060
rect 9294 8032 9295 8043
rect 9294 7964 9295 7975
rect 9303 7914 9304 8094
rect 9305 8066 9306 8100
rect 9667 8092 9668 8126
rect 9812 8100 9813 8111
rect 9656 8058 9657 8069
rect 9823 8066 9824 8100
rect 9979 8092 9980 8126
rect 10124 8100 10125 8111
rect 9968 8058 9969 8069
rect 10135 8066 10136 8100
rect 10291 8092 10292 8126
rect 10436 8100 10437 8111
rect 10280 8058 10281 8069
rect 10447 8066 10448 8100
rect 10603 8092 10604 8126
rect 10748 8100 10749 8111
rect 10592 8058 10593 8069
rect 10759 8066 10760 8100
rect 9305 7998 9306 8032
rect 9667 8024 9668 8058
rect 9812 8032 9813 8043
rect 9656 7990 9657 8001
rect 9823 7998 9824 8032
rect 9979 8024 9980 8058
rect 10124 8032 10125 8043
rect 9968 7990 9969 8001
rect 10135 7998 10136 8032
rect 10291 8024 10292 8058
rect 10436 8032 10437 8043
rect 10280 7990 10281 8001
rect 10447 7998 10448 8032
rect 10603 8024 10604 8058
rect 10748 8032 10749 8043
rect 10592 7990 10593 8001
rect 10759 7998 10760 8032
rect 9305 7930 9306 7964
rect 9667 7956 9668 7990
rect 9812 7964 9813 7975
rect 9656 7922 9657 7933
rect 9823 7930 9824 7964
rect 9979 7956 9980 7990
rect 10124 7964 10125 7975
rect 9968 7922 9969 7933
rect 10135 7930 10136 7964
rect 10291 7956 10292 7990
rect 10436 7964 10437 7975
rect 10280 7922 10281 7933
rect 10447 7930 10448 7964
rect 10603 7956 10604 7990
rect 10748 7964 10749 7975
rect 10592 7922 10593 7933
rect 10759 7930 10760 7964
rect 9667 7888 9668 7922
rect 9979 7888 9980 7922
rect 10291 7888 10292 7922
rect 10603 7888 10604 7922
rect 8202 7716 8203 7727
rect 8213 7682 8214 7716
rect 8358 7710 8359 7721
rect 8514 7716 8515 7727
rect 8369 7676 8370 7710
rect 8525 7682 8526 7716
rect 8670 7710 8671 7721
rect 8826 7716 8827 7727
rect 8681 7676 8682 7710
rect 8837 7682 8838 7716
rect 8982 7710 8983 7721
rect 9138 7716 9139 7727
rect 8993 7676 8994 7710
rect 9149 7682 9150 7716
rect 9628 7702 9629 7713
rect 9940 7702 9941 7713
rect 10252 7702 10253 7713
rect 10592 7702 10593 7713
rect 9639 7668 9640 7702
rect 9951 7668 9952 7702
rect 10263 7668 10264 7702
rect 10603 7668 10604 7702
rect 8202 7648 8203 7659
rect 8213 7614 8214 7648
rect 8358 7642 8359 7653
rect 8514 7648 8515 7659
rect 8369 7608 8370 7642
rect 8525 7614 8526 7648
rect 8670 7642 8671 7653
rect 8826 7648 8827 7659
rect 8681 7608 8682 7642
rect 8837 7614 8838 7648
rect 8982 7642 8983 7653
rect 9138 7648 9139 7659
rect 8993 7608 8994 7642
rect 9149 7614 9150 7648
rect 9628 7634 9629 7645
rect 9784 7642 9785 7653
rect 9639 7600 9640 7634
rect 9795 7608 9796 7642
rect 9940 7634 9941 7645
rect 10096 7642 10097 7653
rect 9951 7600 9952 7634
rect 10107 7608 10108 7642
rect 10252 7634 10253 7645
rect 10408 7642 10409 7653
rect 10263 7600 10264 7634
rect 10419 7608 10420 7642
rect 10592 7634 10593 7645
rect 10603 7600 10604 7634
rect 8071 7528 9345 7578
rect 9479 7528 10799 7578
rect 8071 7454 10837 7456
rect 8289 7146 8489 7196
rect 8575 7146 8775 7196
rect 8787 7146 10391 7196
rect 8339 7100 8340 7145
rect 8724 7134 8725 7145
rect 9092 7134 9093 7145
rect 9404 7134 9405 7145
rect 9716 7134 9717 7145
rect 10028 7134 10029 7145
rect 10340 7134 10341 7145
rect 8735 7100 8736 7134
rect 8936 7092 8937 7103
rect 9103 7100 9104 7134
rect 9248 7092 9249 7103
rect 9415 7100 9416 7134
rect 9560 7092 9561 7103
rect 9727 7100 9728 7134
rect 9872 7092 9873 7103
rect 10039 7100 10040 7134
rect 10184 7092 10185 7103
rect 10351 7100 10352 7134
rect 8071 7016 8169 7066
rect 8339 7026 8340 7071
rect 8724 7066 8725 7077
rect 8735 7032 8736 7066
rect 8947 7058 8948 7092
rect 9092 7066 9093 7077
rect 8936 7024 8937 7035
rect 9103 7032 9104 7066
rect 9259 7058 9260 7092
rect 9404 7066 9405 7077
rect 9248 7024 9249 7035
rect 9415 7032 9416 7066
rect 9571 7058 9572 7092
rect 9716 7066 9717 7077
rect 9560 7024 9561 7035
rect 9727 7032 9728 7066
rect 9883 7058 9884 7092
rect 10028 7066 10029 7077
rect 9872 7024 9873 7035
rect 10039 7032 10040 7066
rect 10195 7058 10196 7092
rect 10340 7066 10341 7077
rect 10184 7024 10185 7035
rect 10351 7032 10352 7066
rect 8724 6998 8725 7009
rect 8339 6952 8340 6997
rect 8735 6964 8736 6998
rect 8947 6990 8948 7024
rect 9092 6998 9093 7009
rect 8936 6956 8937 6967
rect 9103 6964 9104 6998
rect 9259 6990 9260 7024
rect 9404 6998 9405 7009
rect 9248 6956 9249 6967
rect 9415 6964 9416 6998
rect 9571 6990 9572 7024
rect 9716 6998 9717 7009
rect 9560 6956 9561 6967
rect 9727 6964 9728 6998
rect 9883 6990 9884 7024
rect 10028 6998 10029 7009
rect 9872 6956 9873 6967
rect 10039 6964 10040 6998
rect 10195 6990 10196 7024
rect 10340 6998 10341 7009
rect 10184 6956 10185 6967
rect 10351 6964 10352 6998
rect 8724 6930 8725 6941
rect 8339 6874 8340 6919
rect 8735 6896 8736 6930
rect 8947 6922 8948 6956
rect 9092 6930 9093 6941
rect 8936 6888 8937 6899
rect 9103 6896 9104 6930
rect 9259 6922 9260 6956
rect 9404 6930 9405 6941
rect 9248 6888 9249 6899
rect 9415 6896 9416 6930
rect 9571 6922 9572 6956
rect 9716 6930 9717 6941
rect 9560 6888 9561 6899
rect 9727 6896 9728 6930
rect 9883 6922 9884 6956
rect 10028 6930 10029 6941
rect 9872 6888 9873 6899
rect 10039 6896 10040 6930
rect 10195 6922 10196 6956
rect 10340 6930 10341 6941
rect 10184 6888 10185 6899
rect 8071 6816 8169 6866
rect 8947 6854 8948 6888
rect 9259 6854 9260 6888
rect 9571 6854 9572 6888
rect 9883 6854 9884 6888
rect 10195 6854 10196 6888
rect 10315 6846 10316 6896
rect 10349 6880 10350 6930
rect 10351 6896 10352 6930
rect 8936 6668 8937 6679
rect 9092 6676 9093 6687
rect 9248 6682 9249 6693
rect 8071 6578 8123 6628
rect 8339 6610 8340 6655
rect 8947 6634 8948 6668
rect 9103 6642 9104 6676
rect 9259 6648 9260 6682
rect 9404 6676 9405 6687
rect 9560 6682 9561 6693
rect 9415 6642 9416 6676
rect 9571 6648 9572 6682
rect 9716 6676 9717 6687
rect 9872 6682 9873 6693
rect 9727 6642 9728 6676
rect 9883 6648 9884 6682
rect 10028 6676 10029 6687
rect 10184 6682 10185 6693
rect 10039 6642 10040 6676
rect 10195 6648 10196 6682
rect 8936 6600 8937 6611
rect 9092 6608 9093 6619
rect 9248 6614 9249 6625
rect 8339 6542 8340 6587
rect 8947 6566 8948 6600
rect 9103 6574 9104 6608
rect 9259 6580 9260 6614
rect 9404 6608 9405 6619
rect 9560 6614 9561 6625
rect 9415 6574 9416 6608
rect 9571 6580 9572 6614
rect 9716 6608 9717 6619
rect 9872 6614 9873 6625
rect 9727 6574 9728 6608
rect 9883 6580 9884 6614
rect 10028 6608 10029 6619
rect 10184 6614 10185 6625
rect 10039 6574 10040 6608
rect 10195 6580 10196 6614
rect 8289 6460 8489 6510
rect 8579 6494 8779 6544
rect 8787 6494 10391 6544
rect 8073 6420 8107 6422
rect 8169 6420 8203 6422
rect 8265 6420 8299 6422
rect 8361 6420 8395 6422
rect 8457 6420 8491 6422
rect 8553 6420 8587 6422
rect 8649 6420 8683 6422
rect 8745 6420 8779 6422
rect 8841 6420 8875 6422
rect 8937 6420 8971 6422
rect 9033 6420 9067 6422
rect 9129 6420 9163 6422
rect 9225 6420 9259 6422
rect 9321 6420 9355 6422
rect 9417 6420 9451 6422
rect 9513 6420 9547 6422
rect 9609 6420 9643 6422
rect 9705 6420 9739 6422
rect 9801 6420 9835 6422
rect 9897 6420 9931 6422
rect 9993 6420 10027 6422
rect 10089 6420 10123 6422
rect 10185 6420 10219 6422
rect 10281 6420 10315 6422
rect 10377 6420 10411 6422
rect 10473 6420 10507 6422
rect 10569 6420 10603 6422
rect 10665 6420 10699 6422
rect 10761 6420 10795 6422
<< nwell >>
rect 70 7344 6652 7795
rect 7401 6799 10893 7301
<< pwell >>
rect 463 6569 519 6579
rect 2635 5816 2853 6026
<< mvpsubdiff >>
rect 7438 7387 10856 7455
<< mvnsubdiff >>
rect 7467 7201 10827 7235
<< locali >>
rect 41 8275 183 8288
rect 41 8190 57 8275
rect 169 8190 183 8275
rect 41 7451 183 8190
rect 6891 8273 7134 8286
rect 6891 8112 6936 8273
rect 7117 8112 7134 8273
rect 6891 7455 7134 8112
rect 3043 7451 7134 7455
rect 41 7435 7134 7451
rect 41 7305 6927 7435
rect 35 6388 121 7179
rect 3043 7022 6927 7305
rect 7110 7322 7134 7435
rect 7110 7201 10829 7322
rect 7110 7022 7134 7201
rect 3043 7005 7134 7022
rect 2907 6693 7134 6838
rect 2907 6388 3220 6693
rect 35 6320 3220 6388
rect 35 6318 505 6320
rect 35 6192 48 6318
rect 286 6192 505 6318
rect 35 6191 505 6192
rect 2951 6253 3220 6320
rect 6116 6388 7134 6693
rect 6116 6253 10860 6388
rect 2951 6191 10860 6253
rect 35 6143 10860 6191
rect 35 5813 689 6143
rect 1006 5813 1393 6029
rect 1778 5813 2165 6029
rect 2550 6015 2937 6029
rect 2550 5829 2648 6015
rect 2840 5829 2937 6015
rect 2550 5813 2937 5829
rect 3322 5813 3709 6029
rect 4094 5813 4481 6029
rect 4866 5813 5253 6029
rect 5638 5813 6025 6029
rect 6410 5813 6797 6029
rect 7182 5813 7569 6029
rect 7954 5813 8341 6029
rect 8726 5813 9113 6029
rect 9498 5813 9885 6029
rect 10656 5813 10837 6029
rect 51 165 234 381
rect 619 165 1006 381
rect 1391 165 1778 381
rect 2163 165 2550 381
rect 2935 165 3322 381
rect 3707 165 4094 381
rect 4479 165 4866 381
rect 5251 165 5638 381
rect 6023 165 6410 381
rect 6795 165 7182 381
rect 7567 165 7954 381
rect 8339 165 8726 381
rect 9111 165 9498 381
rect 9883 165 10270 381
rect 10655 165 10835 381
<< viali >>
rect 57 8190 169 8275
rect 6936 8112 7117 8273
rect 9224 7854 9270 8060
rect 7604 7754 7807 7801
rect 9459 7754 9796 7801
rect 10785 7683 10819 7879
rect 6927 7022 7110 7435
rect 7870 6775 8128 6834
rect 48 6192 286 6318
rect 505 6191 2951 6320
rect 3220 6253 6116 6693
rect 8439 6684 8506 6878
rect 8650 6720 8853 6767
rect 10270 6735 10316 6896
rect 2648 5829 2840 6015
rect 10202 5598 10340 6030
<< metal1 >>
rect 40 8275 7133 8286
rect 40 8190 57 8275
rect 169 8273 7133 8275
rect 169 8269 6936 8273
rect 624 8260 6936 8269
rect 624 8201 1026 8260
rect 169 8193 1026 8201
rect 7117 8209 7133 8273
rect 7284 8252 10841 8278
rect 169 8190 6936 8193
rect 40 8179 6936 8190
rect 218 8110 376 8127
rect 218 8038 436 8110
rect 709 8082 719 8144
rect 801 8129 818 8144
rect 801 8085 2498 8129
rect 2829 8085 2990 8129
rect 801 8082 818 8085
rect 218 8024 282 8038
rect 218 7641 313 8024
rect 375 7641 436 8038
rect 521 7788 567 8040
rect 627 7892 2821 8028
rect 502 7653 2537 7788
rect 218 7568 436 7641
rect 521 7597 567 7653
rect 709 7597 719 7606
rect 218 7554 375 7568
rect 218 7501 282 7554
rect 521 7553 719 7597
rect 709 7544 719 7553
rect 801 7597 818 7606
rect 2866 7597 2944 8085
rect 2993 7658 3300 7804
rect 801 7556 2990 7597
rect 801 7553 2922 7556
rect 801 7544 818 7553
rect 3360 7501 3433 8122
rect 3699 8082 3959 8128
rect 3486 7636 3556 8035
rect 218 7453 3433 7501
rect 218 7248 282 7453
rect 3497 7344 3556 7636
rect 185 7121 282 7248
rect 2382 7274 3556 7344
rect 3699 7642 3781 8082
rect 4283 8081 5747 8125
rect 6083 8081 6237 8125
rect 6910 8112 6936 8179
rect 7117 8112 7134 8209
rect 7284 8153 7318 8252
rect 10802 8153 10841 8252
rect 7284 8125 10841 8153
rect 3988 7805 4025 8041
rect 4109 7872 6071 8033
rect 3966 7645 5802 7805
rect 3699 7600 3773 7642
rect 3699 7554 3958 7600
rect 3988 7597 4025 7645
rect 6126 7597 6188 8081
rect 6249 7884 6537 8029
rect 6249 7690 6262 7884
rect 3699 7501 3773 7554
rect 3988 7553 6239 7597
rect 6612 7501 6674 8112
rect 3699 7453 6674 7501
rect 185 6969 263 7121
rect 2382 7074 2452 7274
rect 3699 7165 3773 7453
rect 2265 7047 2275 7074
rect 185 6573 282 6969
rect 25 6318 301 6326
rect 25 6192 48 6318
rect 286 6192 301 6318
rect 25 6185 301 6192
rect 25 5348 133 6185
rect 345 5944 399 7033
rect 781 7003 2275 7047
rect 2351 7047 2452 7074
rect 2767 7074 3773 7165
rect 2351 7003 2738 7047
rect 463 6745 634 6972
rect 2382 6952 2452 7003
rect 721 6815 2452 6952
rect 463 6579 2560 6745
rect 463 6569 634 6579
rect 505 6326 634 6569
rect 2629 6533 2693 7003
rect 2767 6949 2842 7074
rect 6752 7065 6823 8044
rect 6910 7435 7134 8112
rect 9218 8060 9276 8072
rect 9218 7854 9224 8060
rect 9270 8051 9276 8060
rect 10128 8051 10138 8053
rect 9270 8001 10138 8051
rect 9270 7854 9276 8001
rect 10128 7999 10138 8001
rect 10290 7999 10300 8053
rect 9218 7842 9276 7854
rect 10779 7879 10825 7891
rect 7592 7801 8339 7807
rect 7592 7754 7604 7801
rect 7807 7754 8339 7801
rect 7592 7748 8339 7754
rect 8519 7801 9808 7807
rect 8519 7754 9459 7801
rect 9796 7754 9808 7801
rect 8519 7748 9808 7754
rect 10779 7728 10785 7879
rect 10819 7728 10825 7879
rect 10743 7674 10753 7728
rect 10905 7674 10915 7728
rect 10779 7671 10825 7674
rect 2756 6573 2842 6949
rect 6407 7036 6825 7065
rect 3167 6819 6174 6842
rect 3167 6693 4331 6819
rect 5278 6693 6174 6819
rect 781 6489 2275 6533
rect 2265 6460 2275 6489
rect 2350 6460 2360 6533
rect 2585 6489 2739 6533
rect 3167 6326 3220 6693
rect 493 6320 3220 6326
rect 493 6191 505 6320
rect 2951 6253 3220 6320
rect 6116 6531 6174 6693
rect 6407 6623 6432 7036
rect 6803 6840 6825 7036
rect 6910 7022 6927 7435
rect 7110 7324 7134 7435
rect 7279 7543 10836 7570
rect 7279 7449 7306 7543
rect 8343 7449 8618 7543
rect 10649 7449 10836 7543
rect 7279 7417 10836 7449
rect 7110 7299 10832 7324
rect 7110 7124 7171 7299
rect 8320 7124 8602 7299
rect 10750 7124 10832 7299
rect 7110 7094 10832 7124
rect 7110 7022 7134 7094
rect 10516 7093 10832 7094
rect 6910 6994 7134 7022
rect 10264 6896 10322 6908
rect 8433 6878 8512 6890
rect 6803 6834 8140 6840
rect 6803 6775 7870 6834
rect 8128 6775 8140 6834
rect 6803 6769 8140 6775
rect 6803 6623 6825 6769
rect 8429 6684 8439 6878
rect 8506 6773 8516 6878
rect 8506 6767 8865 6773
rect 8506 6720 8650 6767
rect 8853 6720 8865 6767
rect 10264 6735 10270 6896
rect 10316 6834 10322 6896
rect 10316 6765 10507 6834
rect 10672 6765 10682 6834
rect 10316 6735 10322 6765
rect 10264 6723 10322 6735
rect 8506 6714 8865 6720
rect 8506 6684 8516 6714
rect 8433 6672 8512 6684
rect 6407 6600 6825 6623
rect 6116 6319 10827 6531
rect 6116 6253 6174 6319
rect 2951 6237 6174 6253
rect 10221 6260 10716 6270
rect 2951 6191 6175 6237
rect 493 6185 6175 6191
rect 10221 6187 10233 6260
rect 10700 6187 10716 6260
rect 10221 6176 10716 6187
rect 10221 6045 10315 6176
rect 10187 6030 10353 6045
rect 2635 6015 2853 6026
rect 2635 5944 2648 6015
rect 345 5890 2648 5944
rect 2635 5829 2648 5890
rect 2840 5829 2853 6015
rect 2635 5816 2853 5829
rect 10187 5598 10202 6030
rect 10340 5598 10353 6030
rect 10187 5582 10353 5598
rect 10805 5348 10867 6079
rect 25 4748 10867 5348
rect 25 4348 133 4748
rect 10805 4348 10867 4748
rect 25 3748 10867 4348
rect 25 3348 133 3748
rect 10805 3348 10867 3748
rect 25 2748 10867 3348
rect 25 2348 133 2748
rect 10805 2348 10867 2748
rect 25 1748 10867 2348
rect 25 1348 133 1748
rect 10805 1348 10867 1748
rect 25 748 10867 1348
rect 25 99 133 748
rect 10805 99 10867 748
rect 25 11 10867 99
<< via1 >>
rect 60 8201 169 8269
rect 169 8201 624 8269
rect 1026 8193 6936 8260
rect 6936 8193 7093 8260
rect 719 8082 801 8144
rect 719 7544 801 7606
rect 7318 8153 10802 8252
rect 2275 7003 2351 7074
rect 10138 7999 10290 8053
rect 8339 7748 8519 7807
rect 10753 7683 10785 7728
rect 10785 7683 10819 7728
rect 10819 7683 10905 7728
rect 10753 7674 10905 7683
rect 4331 6693 5278 6819
rect 2275 6460 2350 6533
rect 4331 6270 5278 6693
rect 6432 6623 6803 7036
rect 7306 7449 8343 7543
rect 8618 7449 10649 7543
rect 7171 7124 8320 7299
rect 8602 7124 10750 7299
rect 8439 6684 8506 6878
rect 10507 6765 10672 6834
rect 10233 6187 10700 6260
<< metal2 >>
rect 985 8286 7132 8287
rect 38 8269 7132 8286
rect 38 8201 60 8269
rect 624 8261 7132 8269
rect 38 8104 77 8201
rect 634 8187 886 8261
rect 7091 8260 7132 8261
rect 7093 8193 7132 8260
rect 634 8104 654 8187
rect 38 8061 654 8104
rect 719 8144 801 8154
rect 719 8072 801 8082
rect 866 8104 886 8187
rect 7091 8104 7132 8193
rect 7284 8252 10841 8278
rect 7284 8153 7318 8252
rect 10802 8153 10841 8252
rect 7284 8125 10841 8153
rect 729 7616 785 8072
rect 866 8060 7132 8104
rect 10138 8056 10290 8066
rect 10138 7986 10290 7996
rect 8339 7807 8519 7817
rect 8339 7738 8519 7748
rect 719 7606 801 7616
rect 719 7534 801 7544
rect 7279 7543 8374 7570
rect 7279 7449 7306 7543
rect 8343 7449 8374 7543
rect 7279 7417 8374 7449
rect 7141 7299 8355 7324
rect 7141 7124 7171 7299
rect 8320 7124 8355 7299
rect 7141 7094 8355 7124
rect 2275 7074 2351 7084
rect 2275 6993 2351 7003
rect 6407 7036 6825 7065
rect 2288 6543 2340 6993
rect 4308 6849 5298 6868
rect 2275 6533 2350 6543
rect 2275 6450 2350 6460
rect 4308 6270 4331 6849
rect 5278 6270 5298 6849
rect 6407 6623 6432 7036
rect 6803 6623 6825 7036
rect 8443 6888 8500 7738
rect 10753 7731 10905 7741
rect 10753 7661 10905 7671
rect 8588 7543 10667 7570
rect 8587 7449 8618 7543
rect 10649 7449 10667 7543
rect 8588 7417 10667 7449
rect 8567 7299 10798 7324
rect 8567 7124 8602 7299
rect 10750 7124 10798 7299
rect 8567 7094 10798 7124
rect 8439 6878 8506 6888
rect 8439 6674 8506 6684
rect 6407 6600 6825 6623
rect 4308 6249 5298 6270
rect 10221 6270 10431 7094
rect 10498 6765 10507 6834
rect 10672 6765 10757 6834
rect 10909 6765 10918 6834
rect 10221 6260 10716 6270
rect 10221 6187 10233 6260
rect 10700 6187 10716 6260
rect 10221 6176 10716 6187
<< via2 >>
rect 77 8201 624 8261
rect 624 8201 634 8261
rect 77 8104 634 8201
rect 886 8260 7091 8261
rect 886 8193 1026 8260
rect 1026 8193 7091 8260
rect 886 8104 7091 8193
rect 7318 8153 10802 8252
rect 10138 8053 10290 8056
rect 10138 7999 10290 8053
rect 10138 7996 10290 7999
rect 7306 7449 8343 7543
rect 4331 6819 5278 6849
rect 4331 6522 5278 6819
rect 6432 6623 6803 7036
rect 10753 7728 10905 7731
rect 10753 7674 10905 7728
rect 10753 7671 10905 7674
rect 8618 7449 10649 7543
rect 10757 6765 10909 6834
<< metal3 >>
rect 38 8261 7126 8283
rect 38 8244 77 8261
rect 634 8244 886 8261
rect 38 8000 73 8244
rect 7091 8104 7126 8261
rect 7284 8252 10841 8278
rect 7284 8153 7318 8252
rect 10802 8153 10841 8252
rect 7284 8125 10841 8153
rect 7073 8000 7126 8104
rect 38 7965 7126 8000
rect 10128 8056 10295 8064
rect 10128 7996 10138 8056
rect 10290 7996 10431 8056
rect 10128 7991 10295 7996
rect 10371 7916 10431 7996
rect 10371 7856 11343 7916
rect 10743 7731 10910 7739
rect 10743 7671 10753 7731
rect 10905 7671 10910 7731
rect 10743 7666 10910 7671
rect 7279 7543 10667 7570
rect 7279 7449 7306 7543
rect 10649 7449 10667 7543
rect 10792 7551 10852 7666
rect 10792 7491 11344 7551
rect 7279 7417 10667 7449
rect 4111 7277 5299 7317
rect 4111 6849 4350 7277
rect 5268 6849 5299 7277
rect 4111 6522 4331 6849
rect 5278 6522 5299 6849
rect 6408 7036 6825 7065
rect 6408 6623 6432 7036
rect 6803 6623 6825 7036
rect 10747 6834 10918 6840
rect 10747 6765 10757 6834
rect 10909 6765 11342 6834
rect 10747 6758 10918 6765
rect 6408 6600 6825 6623
rect 4111 6494 5299 6522
rect 4111 6251 4307 6494
<< via3 >>
rect 73 8104 77 8244
rect 77 8104 634 8244
rect 634 8104 886 8244
rect 886 8104 7073 8244
rect 7318 8153 10802 8252
rect 73 8000 7073 8104
rect 7306 7449 8343 7543
rect 8343 7449 8618 7543
rect 8618 7449 10649 7543
rect 4350 6849 5268 7277
rect 4350 6558 5268 6849
rect 6432 6623 6803 7036
<< metal4 >>
rect 38 8244 7126 8283
rect 38 8000 73 8244
rect 7073 8000 7126 8244
rect 38 7965 7126 8000
rect 7241 8252 11180 8291
rect 7241 8153 7318 8252
rect 10802 8153 11180 8252
rect 7241 7962 11180 8153
rect 10843 7755 11178 7774
rect 38 7543 10667 7655
rect 38 7449 7306 7543
rect 10649 7449 10667 7543
rect 38 7277 10667 7449
rect 38 7255 4350 7277
rect 3817 6558 4350 7255
rect 5268 7255 10667 7277
rect 5268 6558 5299 7255
rect 10843 7074 10879 7755
rect 6386 7036 10879 7074
rect 6386 6623 6432 7036
rect 6803 6623 10879 7036
rect 6386 6615 10879 6623
rect 11146 6615 11178 7755
rect 6386 6591 11178 6615
rect 3817 6522 5299 6558
rect 3817 51 4011 6522
rect 4101 51 4793 6251
<< via4 >>
rect 4350 6558 5268 7247
rect 10879 6615 11146 7755
<< metal5 >>
rect 10851 7755 11171 7779
rect 4313 7247 5299 7317
rect 4313 6558 4350 7247
rect 5268 6558 5299 7247
rect 4313 6494 5299 6558
rect 4507 6135 5299 6494
rect 10851 6615 10879 7755
rect 11146 6615 11171 7755
rect 10851 6242 11171 6615
use sky130_fd_pr__cap_mim_m3_1_WRT4AW  sky130_fd_pr__cap_mim_m3_1_WRT4AW_0
timestamp 1606502073
transform -1 0 7027 0 1 3151
box -3136 -3100 3136 3100
use sky130_fd_pr__cap_mim_m3_2_W5U4AW  sky130_fd_pr__cap_mim_m3_2_W5U4AW_0
timestamp 1606502073
transform 1 0 7970 0 1 3151
box -3179 -3101 3201 3101
use sky130_fd_pr__nfet_g5v0d10v5_PKVMTM  sky130_fd_pr__nfet_g5v0d10v5_PKVMTM_0
timestamp 1606063140
transform 1 0 2660 0 1 6770
box -308 -458 308 458
use sky130_fd_pr__nfet_g5v0d10v5_TGFUGS  sky130_fd_pr__nfet_g5v0d10v5_TGFUGS_0
timestamp 1606063140
transform 1 0 1515 0 1 6769
box -962 -458 962 458
use sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC  sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_1
timestamp 1605994897
transform -1 0 371 0 1 6769
box -308 -458 308 458
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_0
timestamp 1606063140
transform 1 0 3392 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_1
timestamp 1606063140
transform 1 0 3878 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_2
timestamp 1606063140
transform 1 0 6644 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_3
timestamp 1606063140
transform 1 0 408 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_YEUEBV  sky130_fd_pr__pfet_g5v0d10v5_YEUEBV_0
timestamp 1606063140
transform 1 0 5018 0 1 7841
box -992 -497 992 497
use sky130_fd_pr__pfet_g5v0d10v5_YUHPBG  sky130_fd_pr__pfet_g5v0d10v5_YUHPBG_0
timestamp 1606063140
transform 1 0 2906 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_YUHPXE  sky130_fd_pr__pfet_g5v0d10v5_YUHPXE_0
timestamp 1606063140
transform 1 0 6158 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ  sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ_0
timestamp 1606063140
transform 1 0 1657 0 1 7841
box -1101 -497 1101 497
use sky130_fd_pr__res_xhigh_po_0p69_S5N9F3  sky130_fd_pr__res_xhigh_po_0p69_S5N9F3_0
timestamp 1606074388
transform 1 0 5446 0 1 3098
box -5446 -3098 5446 3098
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1681267127
transform 1 0 8523 0 1 6404
box -66 -42 1986 896
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_1
timestamp 1681267127
transform 1 0 7477 0 1 7438
box -66 -42 1986 896
use sky130_fd_sc_hvl__fill_4  sky130_fd_sc_hvl__fill_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1681267127
transform 1 0 10443 0 1 6404
box -66 -42 450 896
use sky130_fd_sc_hvl__inv_8  sky130_fd_sc_hvl__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1681267127
transform 1 0 9397 0 1 7438
box -66 -42 1506 896
use sky130_fd_sc_hvl__schmittbuf_1  sky130_fd_sc_hvl__schmittbuf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1681267127
transform 1 0 7467 0 1 6404
box -66 -42 1122 896
<< labels >>
flabel metal4 s 38 7965 73 8283 0 FreeSans 320 0 0 0 vdd3v3
port 0 nsew
flabel metal4 s 38 7255 232 7655 0 FreeSans 320 0 0 0 vss
port 2 nsew
flabel metal4 s 10974 7962 11180 8291 0 FreeSans 320 0 0 0 vdd1v8
port 1 nsew
flabel metal3 11189 7491 11344 7551 0 FreeSans 320 0 0 0 por_l
port 4 nsew
flabel metal3 11188 7856 11343 7916 0 FreeSans 320 0 0 0 porb_l
port 5 nsew
flabel metal3 10969 6765 11342 6834 0 FreeSans 320 0 0 0 porb_h
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 11344 8338
<< end >>

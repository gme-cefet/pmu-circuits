* NGSPICE file created from ldo.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_lvt_5VYM7K a_n66_n598# a_n124_n510# a_66_n510# VSUBS
X0 a_66_n510# a_n66_n598# a_n124_n510# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
.ends

.subckt sky130_fd_pr__pfet_01v8_TRB9BZ a_n389_n186# w_n483_n189# a_n447_n89# a_389_n89#
+ VSUBS
X0 a_389_n89# a_n389_n186# a_n447_n89# w_n483_n189# sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
C0 a_n389_n186# VSUBS 1.7f
C1 w_n483_n189# VSUBS 1.1f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_8D4JM4 a_n127_n704# w_n221_n707# a_n185_n607#
+ a_127_n607# VSUBS
X0 a_127_n607# a_n127_n704# a_n185_n607# w_n221_n707# sky130_fd_pr__pfet_01v8_lvt ad=1.76 pd=12.7 as=1.76 ps=12.7 w=6.07 l=1.27
C0 w_n221_n707# VSUBS 1.87f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_4FSB7X c1_n546_n1500# m3_n586_n1540# VSUBS
X0 c1_n546_n1500# m3_n586_n1540# sky130_fd_pr__cap_mim_m3_1 l=15 w=4
C0 c1_n546_n1500# m3_n586_n1540# 6.48f
C1 m3_n586_n1540# VSUBS 3.47f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_EFQJD4 a_n95_n517# a_37_n517# a_n37_n614# w_n233_n736#
+ VSUBS
X0 a_37_n517# a_n37_n614# a_n95_n517# w_n233_n736# sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.9 as=1.5 ps=10.9 w=5.17 l=0.37
C0 w_n233_n736# VSUBS 2.92f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_W6ELF5 a_n143_n1235# a_n201_109# a_143_n1147#
+ a_143_109# a_n143_21# a_n201_n1147# a_n303_n1321#
X0 a_143_n1147# a_n143_n1235# a_n201_n1147# a_n303_n1321# sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=5.19 l=1.43
X1 a_143_109# a_n143_21# a_n201_109# a_n303_n1321# sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=5.19 l=1.43
.ends

.subckt ldo Iref VB VS DD OUT SS
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_0 Iref Iref SS SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_1 SS SS SS SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_2 Iref SS m1_9175_n5154# SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_3 Iref SS m1_9116_n8088# SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_5 Iref SS Iref SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_4 Iref SS m1_9116_n8088# SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_6 Iref m1_9116_n8088# SS SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__pfet_01v8_TRB9BZ_0 DD DD DD DD SS sky130_fd_pr__pfet_01v8_TRB9BZ
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_7 Iref m1_9116_n8088# SS SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_8 SS SS SS SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__pfet_01v8_TRB9BZ_2 m1_9175_n5154# DD DD m1_8616_n5605# SS sky130_fd_pr__pfet_01v8_TRB9BZ
Xsky130_fd_pr__pfet_01v8_TRB9BZ_1 DD DD DD DD SS sky130_fd_pr__pfet_01v8_TRB9BZ
Xsky130_fd_pr__nfet_01v8_lvt_5VYM7K_9 Iref m1_9175_n5154# SS SS sky130_fd_pr__nfet_01v8_lvt_5VYM7K
Xsky130_fd_pr__pfet_01v8_TRB9BZ_3 m1_9175_n5154# DD DD m1_9175_n5154# SS sky130_fd_pr__pfet_01v8_TRB9BZ
Xsky130_fd_pr__pfet_01v8_TRB9BZ_4 m1_9175_n5154# DD DD m1_9175_n5154# SS sky130_fd_pr__pfet_01v8_TRB9BZ
Xsky130_fd_pr__pfet_01v8_TRB9BZ_5 m1_9175_n5154# DD DD m1_8616_n5605# SS sky130_fd_pr__pfet_01v8_TRB9BZ
Xsky130_fd_pr__pfet_01v8_lvt_8D4JM4_0 VS OUT OUT m1_9116_n8088# SS sky130_fd_pr__pfet_01v8_lvt_8D4JM4
Xsky130_fd_pr__pfet_01v8_lvt_8D4JM4_1 VS OUT OUT m1_9116_n8088# SS sky130_fd_pr__pfet_01v8_lvt_8D4JM4
Xsky130_fd_pr__cap_mim_m3_1_4FSB7X_0 m1_8616_n5605# OUT SS sky130_fd_pr__cap_mim_m3_1_4FSB7X
Xsky130_fd_pr__pfet_01v8_lvt_EFQJD4_0 DD OUT m1_8616_n5605# DD SS sky130_fd_pr__pfet_01v8_lvt_EFQJD4
Xsky130_fd_pr__nfet_01v8_lvt_W6ELF5_0 VB m1_8616_n5605# m1_9116_n8088# m1_9116_n8088#
+ VB m1_8616_n5605# SS sky130_fd_pr__nfet_01v8_lvt_W6ELF5
X0 m1_9116_n8088# VB.t0 m1_8616_n5605# SS sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=0 l=0
X1 SS Iref.t8 m1_9116_n8088# SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=0 l=0
X2 m1_9116_n8088# Iref.t6 SS SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=0 l=0
X3 DD.t3 DD.t0 DD.t2 DD.t1 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0 l=0
X4 SS Iref.t9 m1_9175_n5154# SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=0 l=0
X5 SS.t7 SS.t4 SS.t6 SS.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=0 l=0
X6 m1_9116_n8088# VS.t0 OUT OUT sky130_fd_pr__pfet_01v8_lvt ad=1.76 pd=12.7 as=1.76 ps=12.7 w=0 l=0
X7 SS Iref.t2 Iref.t3 SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=0 l=0
X8 m1_9116_n8088# Iref.t5 SS SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=0 l=0
X9 SS Iref.t7 m1_9116_n8088# SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=0 l=0
X10 m1_9116_n8088# VS.t1 OUT OUT sky130_fd_pr__pfet_01v8_lvt ad=1.76 pd=12.7 as=1.76 ps=12.7 w=0 l=0
X11 m1_9116_n8088# VB.t1 m1_8616_n5605# SS sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=0 l=0
X12 DD.t7 DD.t4 DD.t6 DD.t5 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0 l=0
X13 SS.t3 SS.t0 SS.t2 SS.t1 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=0 l=0
X14 m1_9175_n5154# Iref.t4 SS SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=0 l=0
X15 Iref.t1 Iref.t0 SS SS sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=0 l=0
R0 Iref.n10 Iref.t4 206.963
R1 Iref.n2 Iref.t9 206.963
R2 Iref.n2 Iref.t7 206.321
R3 Iref.n4 Iref.t8 206.321
R4 Iref.n6 Iref.t2 206.321
R5 Iref.n10 Iref.t5 206.321
R6 Iref.n11 Iref.t6 206.321
R7 Iref.n12 Iref.t0 206.321
R8 Iref.t7 Iref.n1 206.317
R9 Iref.t8 Iref.n3 206.317
R10 Iref.t2 Iref.n5 206.317
R11 Iref.t5 Iref.n9 206.317
R12 Iref.t6 Iref.n8 206.317
R13 Iref.t0 Iref.n7 206.317
R14 Iref.n0 Iref.t1 3.41293
R15 Iref.n0 Iref.t3 3.41293
R16 Iref.n12 Iref.n11 0.642396
R17 Iref.n11 Iref.n10 0.642396
R18 Iref.n4 Iref.n2 0.642396
R19 Iref.n6 Iref.n4 0.642396
R20 Iref.n13 Iref.n12 0.237335
R21 Iref.n13 Iref.n6 0.235494
R22 Iref Iref.n13 0.20576
R23 Iref Iref.n0 0.184094
R24 SS.n19 SS.n18 4862.2
R25 SS.n8 SS.n6 1303.68
R26 SS.n21 SS.n17 774.62
R27 SS.n10 SS.n1 770.619
R28 SS.n24 SS.t1 623.03
R29 SS.n1 SS.n0 610.112
R30 SS.n25 SS.n23 604.529
R31 SS.n17 SS.n14 380.226
R32 SS.n33 SS.n29 340.584
R33 SS.n20 SS.n19 293.863
R34 SS.n27 SS.n21 280.995
R35 SS.n35 SS.n28 270.781
R36 SS.n31 SS.n30 270.476
R37 SS.n9 SS.n4 246.601
R38 SS.n36 SS.n35 227.38
R39 SS.n12 SS.t3 220.899
R40 SS.n30 SS.t0 220.834
R41 SS.n37 SS.t6 220.522
R42 SS.n37 SS.t4 206.317
R43 SS.n43 SS.n42 119.424
R44 SS.n45 SS.n44 102.663
R45 SS.n9 SS.t5 88.811
R46 SS.n28 SS.n27 72.8795
R47 SS.t5 SS.n5 64.6683
R48 SS.n41 SS.n40 56.9082
R49 SS.n27 SS.n26 22.3606
R50 SS.n28 SS.n12 17.6395
R51 SS.n45 SS.n37 17.6395
R52 SS.n22 SS.t2 3.47896
R53 SS.n43 SS.t7 3.41269
R54 SS SS.n36 2.09505
R55 SS.n36 SS.n11 1.88285
R56 SS.n44 SS.n43 1.38918
R57 SS SS.n45 0.756864
R58 SS.n26 SS.n22 0.126275
R59 SS.n26 SS.n25 0.100882
R60 SS.n11 SS.n10 0.0360926
R61 SS.n10 SS.n9 0.0360926
R62 SS.n8 SS.n7 0.0360926
R63 SS.n9 SS.n8 0.0360926
R64 SS.n3 SS.n2 0.00609809
R65 SS.n4 SS.n3 0.00609809
R66 SS.n39 SS.n38 0.00609809
R67 SS.n40 SS.n39 0.00609809
R68 SS.n17 SS.n16 0.00100268
R69 SS.n25 SS.n24 0.00051152
R70 SS.n44 SS.n41 0.00051152
R71 SS.n14 SS.n13 0.000510263
R72 SS.n35 SS.n34 0.000503106
R73 SS.n34 SS.n33 0.000503106
R74 SS.n33 SS.n32 0.000503106
R75 SS.n32 SS.n31 0.000503106
R76 SS.n16 SS.n15 0.000502681
R77 SS.n21 SS.n20 0.000501887
R78 DD.n3 DD.n2 459.671
R79 DD.n22 DD.n16 282.247
R80 DD.n9 DD.n8 254.948
R81 DD.n0 DD.t5 232.912
R82 DD.n7 DD.t1 213.075
R83 DD.n23 DD.n14 209.695
R84 DD.n12 DD.n11 186.632
R85 DD.n10 DD.n9 80.7111
R86 DD.n11 DD.n10 78.8202
R87 DD.n25 DD.n23 63.0245
R88 DD.n2 DD.t3 60.0995
R89 DD.n24 DD.t7 60.0995
R90 DD.n25 DD.n24 53.4946
R91 DD.n9 DD.t2 48.3828
R92 DD.n11 DD.t6 45.276
R93 DD.n23 DD.n22 10.8113
R94 DD.n1 DD.t4 9.47999
R95 DD.n8 DD.t0 9.47999
R96 DD.n26 DD.n25 8.40959
R97 DD.n27 DD.n12 8.10924
R98 DD.n27 DD.n26 5.40633
R99 DD.n12 DD.n1 0.840904
R100 DD DD.n27 0.196382
R101 DD.n14 DD.n13 0.025954
R102 DD.n16 DD.n15 0.025954
R103 DD.n8 DD.n7 0.00450849
R104 DD.n1 DD.n0 0.00450849
R105 DD.n18 DD.n17 0.00414317
R106 DD.n22 DD.n21 0.00414317
R107 DD.n20 DD.n19 0.00397678
R108 DD.n21 DD.n20 0.00355895
R109 DD.n19 DD.n18 0.00348454
R110 DD.n10 DD.n6 0.00193193
R111 DD.n6 DD.n5 0.00193193
R112 DD.n5 DD.n4 0.00193193
R113 DD.n4 DD.n3 0.00193193
R114 VS.n0 VS.t1 147.147
R115 VS.n0 VS.t0 63.6678
R116 VS VS.n0 44.4531
R117 OUT.n7 OUT.n6 261.185
R118 OUT.n2 OUT.n1 229.173
R119 OUT.n10 OUT.n9 74.0415
R120 OUT.n10 OUT.n4 72.1843
R121 OUT.n18 OUT.n10 1.01576
R122 OUT OUT.n18 0.334188
R123 OUT.n4 OUT.n3 0.0153511
R124 OUT.n3 OUT.n2 0.014836
R125 OUT.n9 OUT.n8 0.0131168
R126 OUT.n8 OUT.n7 0.012684
R127 OUT.n18 OUT.n17 0.00718396
R128 OUT.n17 OUT.n16 0.0069195
R129 OUT.n16 OUT.n15 0.00641981
R130 OUT.n17 OUT.n12 0.00449474
R131 OUT.n6 OUT.n5 0.00432563
R132 OUT.n1 OUT.n0 0.00432563
R133 OUT.n12 OUT.n11 0.00399493
R134 OUT.n14 OUT.n13 0.00345991
R135 OUT.n15 OUT.n14 0.00345991
R136 VB.n0 VB.t0 49.9518
R137 VB.n0 VB.t1 48.1905
R138 VB VB.n0 2.76135
C0 OUT m1_8616_n5605# 1.02f
C1 VS OUT 1.62f
C2 m1_8616_n5605# m1_9175_n5154# 1.57f
C3 m1_9116_n8088# OUT 1.41f
C4 m1_9116_n8088# m1_9175_n5154# 1.33f
C5 OUT VB 1.46f
C6 VB m1_9175_n5154# 1.24f
C7 m1_9116_n8088# VB 3.13f
C8 DD m1_8616_n5605# 1.26f
C9 DD m1_9175_n5154# 3.18f
C10 Iref SS 6.7f
C11 DD SS 20.7f
C12 VB.n0 SS 1.72f
C13 OUT.n18 SS 4.73f
C14 m1_8616_n5605# SS 4.94f
C15 VB SS 4.87f
C16 VS SS 1.28f
C17 OUT SS 14.6f
C18 m1_9116_n8088# SS 6.66f
C19 m1_9175_n5154# SS 6.36f
.ends


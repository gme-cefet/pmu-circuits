magic
tech sky130A
magscale 1 2
timestamp 1697399585
<< nwell >>
rect -195 -195 195 195
<< pwell >>
rect -333 195 333 333
rect -333 -195 -195 195
rect 195 -195 333 195
rect -333 -333 333 -195
<< psubdiff >>
rect -297 263 -201 297
rect 201 263 297 297
rect -297 201 -263 263
rect 263 201 297 263
rect -297 -263 -263 -201
rect 263 -263 297 -201
rect -297 -297 -201 -263
rect 201 -297 297 -263
<< nsubdiff >>
rect -159 147 159 159
rect -159 113 -51 147
rect 51 113 159 147
rect -159 101 159 113
rect -159 51 -101 101
rect -159 -51 -147 51
rect -113 -51 -101 51
rect 101 51 159 101
rect -159 -101 -101 -51
rect 101 -51 113 51
rect 147 -51 159 51
rect 101 -101 159 -51
rect -159 -113 159 -101
rect -159 -147 -51 -113
rect 51 -147 159 -113
rect -159 -159 159 -147
<< psubdiffcont >>
rect -201 263 201 297
rect -297 -201 -263 201
rect 263 -201 297 201
rect -201 -297 201 -263
<< nsubdiffcont >>
rect -51 113 51 147
rect -147 -51 -113 51
rect 113 -51 147 51
rect -51 -147 51 -113
<< pdiodelvt >>
rect -45 33 45 45
rect -45 -33 -33 33
rect 33 -33 45 33
rect -45 -45 45 -33
<< pdiodelvtc >>
rect -33 -33 33 33
<< locali >>
rect -297 263 -201 297
rect 201 263 297 297
rect -297 201 -263 263
rect 263 201 297 263
rect -147 113 -51 147
rect 51 113 147 147
rect -147 51 -113 113
rect 113 51 147 113
rect -49 -33 -33 33
rect 33 -33 49 33
rect -147 -113 -113 -51
rect 113 -113 147 -51
rect -147 -147 -51 -113
rect 51 -147 147 -113
rect -297 -263 -263 -201
rect 263 -263 297 -201
rect -297 -297 -201 -263
rect 201 -297 297 -263
<< viali >>
rect -33 -33 33 33
<< metal1 >>
rect -45 33 45 39
rect -45 -33 -33 33
rect 33 -33 45 33
rect -45 -39 45 -33
<< properties >>
string FIXED_BBOX -130 -130 130 130
string gencell sky130_fd_pr__diode_pd2nw_05v5_lvt
string library sky130
string parameters w 0.45 l 0.45 area 202.5m peri 1.8 nx 1 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 0 compatible {sky130_fd_pr__diode_pd2nw_05v5 sky130_fd_pr__diode_pd2nw_05v5_lvt  sky130_fd_pr__diode_pd2nw_05v5_hvt sky130_fd_pr__diode_pd2nw_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

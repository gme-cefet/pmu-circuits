magic
tech sky130A
magscale 1 2
timestamp 1697059543
<< nwell >>
rect -1334 -3224 33 -1036
rect 297 -2846 911 -1060
rect 1177 -3811 1669 -1065
<< pmos >>
rect -1082 -2108 -608 -1232
rect 1373 -1684 1473 -1284
rect 1373 -2320 1473 -1920
rect 1373 -2956 1473 -2556
rect 1373 -3592 1473 -3192
<< pmoslvt >>
rect -316 -2034 -216 -1234
rect -896 -3028 -210 -2474
rect 516 -2650 692 -1256
<< pdiff >>
rect -1082 -1186 -608 -1174
rect -1082 -1220 -1070 -1186
rect -620 -1220 -608 -1186
rect -1082 -1232 -608 -1220
rect -316 -1188 -216 -1176
rect -316 -1222 -304 -1188
rect -228 -1222 -216 -1188
rect -316 -1234 -216 -1222
rect -316 -2046 -216 -2034
rect -316 -2080 -304 -2046
rect -228 -2080 -216 -2046
rect -316 -2092 -216 -2080
rect -1082 -2120 -608 -2108
rect -1082 -2154 -1070 -2120
rect -620 -2154 -608 -2120
rect -1082 -2166 -608 -2154
rect -896 -2428 -210 -2416
rect -896 -2462 -884 -2428
rect -222 -2462 -210 -2428
rect -896 -2474 -210 -2462
rect -896 -3040 -210 -3028
rect -896 -3074 -884 -3040
rect -222 -3074 -210 -3040
rect -896 -3086 -210 -3074
rect 516 -1210 692 -1198
rect 516 -1244 528 -1210
rect 680 -1244 692 -1210
rect 516 -1256 692 -1244
rect 516 -2662 692 -2650
rect 516 -2696 528 -2662
rect 680 -2696 692 -2662
rect 516 -2708 692 -2696
rect 1315 -1296 1373 -1284
rect 1315 -1672 1327 -1296
rect 1361 -1672 1373 -1296
rect 1315 -1684 1373 -1672
rect 1473 -1296 1531 -1284
rect 1473 -1672 1485 -1296
rect 1519 -1672 1531 -1296
rect 1473 -1684 1531 -1672
rect 1315 -1932 1373 -1920
rect 1315 -2308 1327 -1932
rect 1361 -2308 1373 -1932
rect 1315 -2320 1373 -2308
rect 1473 -1932 1531 -1920
rect 1473 -2308 1485 -1932
rect 1519 -2308 1531 -1932
rect 1473 -2320 1531 -2308
rect 1315 -2568 1373 -2556
rect 1315 -2944 1327 -2568
rect 1361 -2944 1373 -2568
rect 1315 -2956 1373 -2944
rect 1473 -2568 1531 -2556
rect 1473 -2944 1485 -2568
rect 1519 -2944 1531 -2568
rect 1473 -2956 1531 -2944
rect 1315 -3204 1373 -3192
rect 1315 -3580 1327 -3204
rect 1361 -3580 1373 -3204
rect 1315 -3592 1373 -3580
rect 1473 -3204 1531 -3192
rect 1473 -3580 1485 -3204
rect 1519 -3580 1531 -3204
rect 1473 -3592 1531 -3580
<< pdiffc >>
rect -1070 -1220 -620 -1186
rect -304 -1222 -228 -1188
rect -304 -2080 -228 -2046
rect -1070 -2154 -620 -2120
rect -884 -2462 -222 -2428
rect -884 -3074 -222 -3040
rect 528 -1244 680 -1210
rect 528 -2696 680 -2662
rect 1327 -1672 1361 -1296
rect 1485 -1672 1519 -1296
rect 1327 -2308 1361 -1932
rect 1485 -2308 1519 -1932
rect 1327 -2944 1361 -2568
rect 1485 -2944 1519 -2568
rect 1327 -3580 1361 -3204
rect 1485 -3580 1519 -3204
<< psubdiff >>
rect -1459 -962 -1435 -845
rect 1653 -962 1677 -845
<< nsubdiff >>
rect -1298 -1106 -1238 -1072
rect -63 -1106 -3 -1072
rect -1298 -1132 -1264 -1106
rect -37 -1132 -3 -1106
rect -1298 -3154 -1264 -3128
rect 333 -1130 429 -1096
rect 779 -1130 875 -1096
rect 333 -1192 367 -1130
rect 841 -1192 875 -1130
rect 333 -2776 367 -2714
rect 841 -2776 875 -2714
rect 333 -2810 429 -2776
rect 779 -2810 875 -2776
rect 1213 -1135 1309 -1101
rect 1537 -1135 1633 -1101
rect 1213 -1197 1247 -1135
rect -37 -3154 -3 -3128
rect -1298 -3188 -1238 -3154
rect -63 -3188 -3 -3154
rect 1599 -1197 1633 -1135
rect 1213 -3741 1247 -3679
rect 1599 -3741 1633 -3679
rect 1213 -3775 1309 -3741
rect 1537 -3775 1633 -3741
<< psubdiffcont >>
rect -1435 -962 1653 -845
<< nsubdiffcont >>
rect -1238 -1106 -63 -1072
rect -1298 -3128 -1264 -1132
rect -37 -3128 -3 -1132
rect 429 -1130 779 -1096
rect 333 -2714 367 -1192
rect 841 -2714 875 -1192
rect 429 -2810 779 -2776
rect 1309 -1135 1537 -1101
rect -1238 -3188 -63 -3154
rect 1213 -3679 1247 -1197
rect 1599 -3679 1633 -1197
rect 1309 -3775 1537 -3741
<< poly >>
rect -1179 -1248 -1082 -1232
rect -1179 -2092 -1163 -1248
rect -1129 -2092 -1082 -1248
rect -1179 -2108 -1082 -2092
rect -608 -1248 -511 -1232
rect -608 -2092 -561 -1248
rect -527 -2092 -511 -1248
rect -413 -1250 -316 -1234
rect -413 -2018 -397 -1250
rect -363 -2018 -316 -1250
rect -413 -2034 -316 -2018
rect -216 -1250 -119 -1234
rect -216 -2018 -169 -1250
rect -135 -2018 -119 -1250
rect -216 -2034 -119 -2018
rect -608 -2108 -511 -2092
rect -993 -2490 -896 -2474
rect -993 -3012 -977 -2490
rect -943 -3012 -896 -2490
rect -993 -3028 -896 -3012
rect -210 -2490 -113 -2474
rect -210 -3012 -163 -2490
rect -129 -3012 -113 -2490
rect -210 -3028 -113 -3012
rect 419 -1272 516 -1256
rect 419 -2634 435 -1272
rect 469 -2634 516 -1272
rect 419 -2650 516 -2634
rect 692 -1272 789 -1256
rect 692 -2634 739 -1272
rect 773 -2634 789 -1272
rect 692 -2650 789 -2634
rect 1373 -1203 1473 -1187
rect 1373 -1237 1389 -1203
rect 1457 -1237 1473 -1203
rect 1373 -1284 1473 -1237
rect 1373 -1731 1473 -1684
rect 1373 -1765 1389 -1731
rect 1457 -1765 1473 -1731
rect 1373 -1781 1473 -1765
rect 1373 -1839 1473 -1823
rect 1373 -1873 1389 -1839
rect 1457 -1873 1473 -1839
rect 1373 -1920 1473 -1873
rect 1373 -2367 1473 -2320
rect 1373 -2401 1389 -2367
rect 1457 -2401 1473 -2367
rect 1373 -2417 1473 -2401
rect 1373 -2475 1473 -2459
rect 1373 -2509 1389 -2475
rect 1457 -2509 1473 -2475
rect 1373 -2556 1473 -2509
rect 1373 -3003 1473 -2956
rect 1373 -3037 1389 -3003
rect 1457 -3037 1473 -3003
rect 1373 -3053 1473 -3037
rect 1373 -3111 1473 -3095
rect 1373 -3145 1389 -3111
rect 1457 -3145 1473 -3111
rect 1373 -3192 1473 -3145
rect 1373 -3639 1473 -3592
rect 1373 -3673 1389 -3639
rect 1457 -3673 1473 -3639
rect 1373 -3689 1473 -3673
<< polycont >>
rect -1163 -2092 -1129 -1248
rect -561 -2092 -527 -1248
rect -397 -2018 -363 -1250
rect -169 -2018 -135 -1250
rect -977 -3012 -943 -2490
rect -163 -3012 -129 -2490
rect 435 -2634 469 -1272
rect 739 -2634 773 -1272
rect 1389 -1237 1457 -1203
rect 1389 -1765 1457 -1731
rect 1389 -1873 1457 -1839
rect 1389 -2401 1457 -2367
rect 1389 -2509 1457 -2475
rect 1389 -3037 1457 -3003
rect 1389 -3145 1457 -3111
rect 1389 -3673 1457 -3639
<< locali >>
rect -1451 -962 -1435 -845
rect 1653 -962 1669 -845
rect -1298 -1078 -1238 -1072
rect -1434 -1106 -1238 -1078
rect -63 -1106 -3 -1072
rect -1434 -1132 -1264 -1106
rect -1434 -2176 -1298 -1132
rect -922 -1186 -749 -1106
rect -1086 -1220 -1070 -1186
rect -620 -1220 -604 -1186
rect -283 -1188 -239 -1106
rect -37 -1132 -3 -1106
rect -320 -1222 -304 -1188
rect -228 -1222 -212 -1188
rect -1163 -1248 -1129 -1232
rect -1163 -2108 -1129 -2092
rect -561 -1248 -527 -1232
rect -397 -1250 -363 -1234
rect -397 -2034 -363 -2018
rect -169 -1250 -135 -1234
rect -169 -2034 -135 -2018
rect -320 -2080 -304 -2046
rect -228 -2080 -212 -2046
rect -561 -2108 -527 -2092
rect -1086 -2154 -1070 -2120
rect -620 -2154 -604 -2120
rect -1009 -2312 -970 -2154
rect -1009 -2353 -106 -2312
rect -1009 -2474 -970 -2353
rect -900 -2462 -884 -2428
rect -222 -2462 -206 -2428
rect -146 -2474 -106 -2353
rect -1009 -2490 -943 -2474
rect -1009 -3012 -977 -2490
rect -1009 -3028 -943 -3012
rect -163 -2490 -106 -2474
rect -129 -3012 -106 -2490
rect -163 -3028 -106 -3012
rect -900 -3074 -884 -3040
rect -222 -3074 -206 -3040
rect -1298 -3154 -1264 -3128
rect 333 -1130 429 -1096
rect 779 -1130 875 -1096
rect 333 -1192 875 -1130
rect 108 -2554 333 -2504
rect 108 -2731 150 -2554
rect 303 -2714 333 -2554
rect 367 -1210 841 -1192
rect 367 -1244 528 -1210
rect 680 -1244 841 -1210
rect 367 -1272 469 -1244
rect 367 -2634 435 -1272
rect 367 -2650 469 -2634
rect 739 -1272 841 -1244
rect 773 -2634 841 -1272
rect 739 -2650 841 -2634
rect 367 -2678 444 -2650
rect 512 -2696 528 -2662
rect 680 -2696 696 -2662
rect 765 -2680 841 -2650
rect 303 -2731 367 -2714
rect 108 -2763 367 -2731
rect 333 -2776 367 -2763
rect 1030 -1222 1053 -962
rect 1124 -1222 1149 -962
rect 1030 -1245 1149 -1222
rect 1213 -1135 1309 -1101
rect 1537 -1135 1633 -1101
rect 1213 -1197 1247 -1135
rect 841 -2776 875 -2714
rect 333 -2810 429 -2776
rect 779 -2810 875 -2776
rect -37 -3154 -3 -3128
rect -1298 -3188 -1238 -3154
rect -63 -3188 -3 -3154
rect 1074 -3283 1213 -3263
rect 1074 -3367 1101 -3283
rect 1202 -3367 1213 -3283
rect 1074 -3385 1213 -3367
rect 1599 -1197 1633 -1135
rect 1373 -1237 1389 -1203
rect 1457 -1237 1473 -1203
rect 1327 -1296 1361 -1280
rect 1327 -1688 1361 -1672
rect 1485 -1296 1599 -1280
rect 1519 -1672 1599 -1296
rect 1485 -1688 1599 -1672
rect 1373 -1765 1389 -1731
rect 1457 -1765 1473 -1731
rect 1373 -1873 1389 -1839
rect 1457 -1873 1473 -1839
rect 1327 -1932 1361 -1916
rect 1327 -2324 1361 -2308
rect 1485 -1932 1599 -1916
rect 1519 -2308 1599 -1932
rect 1485 -2324 1599 -2308
rect 1373 -2401 1389 -2367
rect 1457 -2401 1473 -2367
rect 1373 -2509 1389 -2475
rect 1457 -2509 1473 -2475
rect 1327 -2568 1361 -2552
rect 1327 -2960 1361 -2944
rect 1485 -2568 1599 -2552
rect 1519 -2944 1599 -2568
rect 1485 -2960 1599 -2944
rect 1373 -3037 1389 -3003
rect 1457 -3037 1473 -3003
rect 1373 -3145 1389 -3111
rect 1457 -3145 1473 -3111
rect 1327 -3204 1361 -3188
rect 1327 -3596 1361 -3580
rect 1485 -3204 1599 -3188
rect 1519 -3580 1599 -3204
rect 1485 -3596 1599 -3580
rect 1373 -3673 1389 -3639
rect 1457 -3673 1473 -3639
rect 1213 -3741 1247 -3679
rect 1599 -3741 1633 -3679
rect 1213 -3775 1309 -3741
rect 1537 -3775 1633 -3741
<< viali >>
rect 1053 -962 1124 -938
rect -1070 -1220 -620 -1186
rect -304 -1222 -228 -1188
rect -1163 -2092 -1129 -1248
rect -561 -2092 -527 -1248
rect -397 -2018 -363 -1250
rect -169 -2018 -135 -1250
rect -304 -2080 -228 -2046
rect -1070 -2154 -620 -2120
rect -884 -2462 -222 -2428
rect -977 -3012 -943 -2490
rect -163 -3012 -129 -2490
rect -884 -3074 -222 -3040
rect 150 -2731 303 -2554
rect 528 -1244 680 -1210
rect 435 -2634 469 -1272
rect 739 -2634 773 -1272
rect 528 -2696 680 -2662
rect 1053 -1222 1124 -962
rect 1101 -3367 1202 -3283
rect 1389 -1237 1457 -1203
rect 1327 -1672 1361 -1296
rect 1485 -1672 1519 -1296
rect 1389 -1765 1457 -1731
rect 1389 -1873 1457 -1839
rect 1327 -2308 1361 -1932
rect 1485 -2308 1519 -1932
rect 1389 -2401 1457 -2367
rect 1389 -2509 1457 -2475
rect 1327 -2944 1361 -2568
rect 1485 -2944 1519 -2568
rect 1389 -3037 1457 -3003
rect 1389 -3145 1457 -3111
rect 1327 -3580 1361 -3204
rect 1485 -3580 1519 -3204
rect 1389 -3673 1457 -3639
<< metal1 >>
rect 1030 -938 1149 -914
rect -1082 -1186 -608 -1180
rect -1082 -1220 -1070 -1186
rect -620 -1220 -608 -1186
rect -1082 -1226 -608 -1220
rect -403 -1188 -129 -1182
rect -403 -1222 -304 -1188
rect -228 -1222 -129 -1188
rect -403 -1228 -129 -1222
rect -1169 -1248 -1123 -1236
rect -1169 -1280 -1163 -1248
rect -1200 -2092 -1163 -1280
rect -1129 -2092 -1123 -1248
rect -1200 -2104 -1123 -2092
rect -567 -1248 -486 -1236
rect -567 -2092 -561 -1248
rect -527 -2092 -486 -1248
rect -403 -1238 -316 -1228
rect -216 -1238 -129 -1228
rect -403 -1250 -357 -1238
rect -403 -2018 -397 -1250
rect -363 -2018 -357 -1250
rect -403 -2030 -357 -2018
rect -175 -1250 -129 -1238
rect 516 -1210 692 -1204
rect 516 -1244 528 -1210
rect 680 -1244 692 -1210
rect 516 -1250 692 -1244
rect 1030 -1222 1053 -938
rect 1124 -1208 1149 -938
rect 1377 -1203 1469 -1197
rect 1377 -1208 1389 -1203
rect 1124 -1222 1389 -1208
rect 1030 -1237 1389 -1222
rect 1457 -1237 1469 -1203
rect 1030 -1240 1469 -1237
rect 1030 -1245 1149 -1240
rect 1377 -1243 1469 -1240
rect -175 -2018 -169 -1250
rect -135 -2018 -129 -1250
rect -175 -2030 -129 -2018
rect 429 -1272 475 -1260
rect -567 -2104 -486 -2092
rect -1200 -2258 -1158 -2104
rect -1082 -2120 -608 -2114
rect -1082 -2154 -1070 -2120
rect -620 -2154 -608 -2120
rect -1082 -2160 -608 -2154
rect -523 -2258 -486 -2104
rect -316 -2046 -216 -2040
rect -316 -2080 -304 -2046
rect -228 -2080 -216 -2046
rect -316 -2258 -216 -2080
rect -1200 -2295 -216 -2258
rect -316 -2422 -216 -2295
rect -896 -2428 -210 -2422
rect -896 -2462 -884 -2428
rect -222 -2462 -210 -2428
rect -896 -2468 -210 -2462
rect -983 -2490 -937 -2478
rect -983 -3012 -977 -2490
rect -943 -3012 -937 -2490
rect -983 -3024 -937 -3012
rect -169 -2490 -123 -2478
rect -169 -3012 -163 -2490
rect -129 -2610 -123 -2490
rect 108 -2554 347 -2504
rect 108 -2610 150 -2554
rect -129 -2731 150 -2610
rect 303 -2731 347 -2554
rect 429 -2634 435 -1272
rect 469 -2634 475 -1272
rect 429 -2646 475 -2634
rect 733 -1272 779 -1260
rect 733 -2634 739 -1272
rect 773 -2634 779 -1272
rect 733 -2646 779 -2634
rect 1066 -1447 1135 -1245
rect 1321 -1296 1367 -1284
rect 1321 -1447 1327 -1296
rect 1066 -1504 1327 -1447
rect 1066 -1788 1135 -1504
rect 1321 -1672 1327 -1504
rect 1361 -1672 1367 -1296
rect 1321 -1684 1367 -1672
rect 1479 -1296 1525 -1284
rect 1479 -1672 1485 -1296
rect 1519 -1672 1525 -1296
rect 1479 -1684 1525 -1672
rect 1377 -1731 1469 -1725
rect 1377 -1765 1389 -1731
rect 1457 -1765 1469 -1731
rect 1377 -1788 1469 -1765
rect 1066 -1820 1469 -1788
rect 1066 -2090 1135 -1820
rect 1377 -1839 1469 -1820
rect 1377 -1873 1389 -1839
rect 1457 -1873 1469 -1839
rect 1377 -1879 1469 -1873
rect 1321 -1932 1367 -1920
rect 1321 -2090 1327 -1932
rect 1066 -2147 1327 -2090
rect 1066 -2423 1135 -2147
rect 1321 -2308 1327 -2147
rect 1361 -2308 1367 -1932
rect 1321 -2320 1367 -2308
rect 1479 -1932 1525 -1920
rect 1479 -2308 1485 -1932
rect 1519 -2308 1525 -1932
rect 1479 -2320 1525 -2308
rect 1377 -2367 1469 -2361
rect 1377 -2401 1389 -2367
rect 1457 -2401 1469 -2367
rect 1377 -2423 1469 -2401
rect 1066 -2455 1469 -2423
rect 516 -2662 692 -2656
rect 516 -2696 528 -2662
rect 680 -2696 692 -2662
rect 516 -2702 692 -2696
rect -129 -2763 347 -2731
rect -129 -3012 -123 -2763
rect 538 -2873 670 -2702
rect 1066 -2733 1135 -2455
rect 1377 -2475 1469 -2455
rect 1377 -2509 1389 -2475
rect 1457 -2509 1469 -2475
rect 1377 -2515 1469 -2509
rect 1321 -2568 1367 -2556
rect 1321 -2733 1327 -2568
rect 1066 -2790 1327 -2733
rect 1066 -2873 1135 -2790
rect 538 -2930 1135 -2873
rect -169 -3024 -123 -3012
rect -896 -3040 -210 -3034
rect -896 -3074 -884 -3040
rect -222 -3074 -210 -3040
rect -896 -3080 -210 -3074
rect -344 -3263 -210 -3080
rect 1066 -3058 1135 -2930
rect 1321 -2944 1327 -2790
rect 1361 -2944 1367 -2568
rect 1321 -2956 1367 -2944
rect 1479 -2568 1525 -2556
rect 1479 -2944 1485 -2568
rect 1519 -2944 1525 -2568
rect 1479 -2956 1525 -2944
rect 1377 -3003 1469 -2997
rect 1377 -3037 1389 -3003
rect 1457 -3037 1469 -3003
rect 1377 -3058 1469 -3037
rect 1066 -3062 1469 -3058
rect 1066 -3090 1752 -3062
rect 1066 -3167 1135 -3090
rect 1321 -3103 1752 -3090
rect 1321 -3111 1469 -3103
rect 1321 -3145 1389 -3111
rect 1457 -3145 1469 -3111
rect 1321 -3151 1469 -3145
rect 1321 -3192 1387 -3151
rect 1321 -3204 1367 -3192
rect -344 -3283 1229 -3263
rect -344 -3367 1101 -3283
rect 1202 -3367 1229 -3283
rect -344 -3385 1229 -3367
rect 1321 -3580 1327 -3204
rect 1361 -3580 1367 -3204
rect 1321 -3592 1367 -3580
rect 1479 -3204 1525 -3192
rect 1479 -3580 1485 -3204
rect 1519 -3580 1525 -3204
rect 1479 -3592 1525 -3580
rect 1377 -3636 1469 -3633
rect 1709 -3636 1752 -3103
rect 1377 -3639 1752 -3636
rect 1377 -3673 1389 -3639
rect 1457 -3673 1752 -3639
rect 1377 -3677 1752 -3673
rect 1377 -3679 1469 -3677
<< labels >>
flabel locali -1422 -1274 -1344 -1196 0 FreeSans 1600 0 0 0 DD
port 0 nsew
flabel locali 540 -952 626 -878 0 FreeSans 1600 0 0 0 SS
port 1 nsew
flabel metal1 552 -3360 638 -3286 0 FreeSans 1600 0 0 0 VREF
port 2 nsew
<< end >>

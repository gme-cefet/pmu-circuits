magic
tech sky130A
magscale 1 2
timestamp 1695321174
<< error_p >>
rect 486 8166 1778 8216
rect 1940 8166 3214 8216
rect 536 8154 537 8165
rect 848 8154 849 8165
rect 1160 8154 1161 8165
rect 1472 8154 1473 8165
rect 1990 8154 1991 8165
rect 2302 8154 2303 8165
rect 2614 8154 2615 8165
rect 2926 8154 2927 8165
rect 22203 8158 23477 8208
rect 23639 8158 24931 8208
rect 525 8120 526 8154
rect 692 8112 693 8123
rect 837 8120 838 8154
rect 1004 8112 1005 8123
rect 1149 8120 1150 8154
rect 1316 8112 1317 8123
rect 1461 8120 1462 8154
rect 1628 8112 1629 8123
rect 1979 8120 1980 8154
rect 2146 8112 2147 8123
rect 2291 8120 2292 8154
rect 2458 8112 2459 8123
rect 2603 8120 2604 8154
rect 2770 8112 2771 8123
rect 2915 8120 2916 8154
rect 22490 8146 22491 8157
rect 22802 8146 22803 8157
rect 23114 8146 23115 8157
rect 23426 8146 23427 8157
rect 23944 8146 23945 8157
rect 24256 8146 24257 8157
rect 24568 8146 24569 8157
rect 24880 8146 24881 8157
rect 3082 8112 3083 8123
rect 536 8086 537 8097
rect 525 8052 526 8086
rect 681 8078 682 8112
rect 848 8086 849 8097
rect 692 8044 693 8055
rect 837 8052 838 8086
rect 993 8078 994 8112
rect 1160 8086 1161 8097
rect 1004 8044 1005 8055
rect 1149 8052 1150 8086
rect 1305 8078 1306 8112
rect 1472 8086 1473 8097
rect 1316 8044 1317 8055
rect 1461 8052 1462 8086
rect 1617 8078 1618 8112
rect 1990 8086 1991 8097
rect 1628 8044 1629 8055
rect 1979 8052 1980 8086
rect 536 8018 537 8029
rect 525 7984 526 8018
rect 681 8010 682 8044
rect 848 8018 849 8029
rect 692 7976 693 7987
rect 837 7984 838 8018
rect 993 8010 994 8044
rect 1160 8018 1161 8029
rect 1004 7976 1005 7987
rect 1149 7984 1150 8018
rect 1305 8010 1306 8044
rect 1472 8018 1473 8029
rect 1316 7976 1317 7987
rect 1461 7984 1462 8018
rect 1617 8010 1618 8044
rect 1628 7976 1629 7987
rect 1979 7984 1980 8018
rect 536 7950 537 7961
rect 525 7916 526 7950
rect 681 7942 682 7976
rect 848 7950 849 7961
rect 692 7908 693 7919
rect 837 7916 838 7950
rect 993 7942 994 7976
rect 1160 7950 1161 7961
rect 1004 7908 1005 7919
rect 1149 7916 1150 7950
rect 1305 7942 1306 7976
rect 1472 7950 1473 7961
rect 1316 7908 1317 7919
rect 1461 7916 1462 7950
rect 1617 7942 1618 7976
rect 1628 7908 1629 7919
rect 1979 7916 1980 7950
rect 681 7874 682 7908
rect 993 7874 994 7908
rect 1305 7874 1306 7908
rect 1617 7874 1618 7908
rect 1981 7900 1982 8080
rect 2135 8078 2136 8112
rect 2302 8086 2303 8097
rect 1990 8018 1991 8029
rect 1990 7950 1991 7961
rect 2015 7866 2016 8046
rect 2146 8044 2147 8055
rect 2291 8052 2292 8086
rect 2447 8078 2448 8112
rect 2614 8086 2615 8097
rect 2458 8044 2459 8055
rect 2603 8052 2604 8086
rect 2759 8078 2760 8112
rect 2926 8086 2927 8097
rect 2770 8044 2771 8055
rect 2915 8052 2916 8086
rect 3071 8078 3072 8112
rect 22334 8104 22335 8115
rect 22501 8112 22502 8146
rect 22646 8104 22647 8115
rect 22813 8112 22814 8146
rect 22958 8104 22959 8115
rect 23125 8112 23126 8146
rect 23270 8104 23271 8115
rect 23437 8112 23438 8146
rect 23788 8104 23789 8115
rect 23955 8112 23956 8146
rect 24100 8104 24101 8115
rect 24267 8112 24268 8146
rect 24412 8104 24413 8115
rect 24579 8112 24580 8146
rect 24724 8104 24725 8115
rect 24891 8112 24892 8146
rect 22345 8070 22346 8104
rect 22490 8078 22491 8089
rect 3082 8044 3083 8055
rect 2135 8010 2136 8044
rect 2302 8018 2303 8029
rect 2146 7976 2147 7987
rect 2291 7984 2292 8018
rect 2447 8010 2448 8044
rect 2614 8018 2615 8029
rect 2458 7976 2459 7987
rect 2603 7984 2604 8018
rect 2759 8010 2760 8044
rect 2926 8018 2927 8029
rect 2770 7976 2771 7987
rect 2915 7984 2916 8018
rect 3071 8010 3072 8044
rect 22334 8036 22335 8047
rect 22501 8044 22502 8078
rect 22657 8070 22658 8104
rect 22802 8078 22803 8089
rect 22646 8036 22647 8047
rect 22813 8044 22814 8078
rect 22969 8070 22970 8104
rect 23114 8078 23115 8089
rect 22958 8036 22959 8047
rect 23125 8044 23126 8078
rect 23281 8070 23282 8104
rect 23426 8078 23427 8089
rect 23270 8036 23271 8047
rect 22345 8002 22346 8036
rect 22490 8010 22491 8021
rect 3082 7976 3083 7987
rect 2135 7942 2136 7976
rect 2302 7950 2303 7961
rect 2146 7908 2147 7919
rect 2291 7916 2292 7950
rect 2447 7942 2448 7976
rect 2614 7950 2615 7961
rect 2458 7908 2459 7919
rect 2603 7916 2604 7950
rect 2759 7942 2760 7976
rect 2926 7950 2927 7961
rect 2770 7908 2771 7919
rect 2915 7916 2916 7950
rect 3071 7942 3072 7976
rect 22334 7968 22335 7979
rect 22501 7976 22502 8010
rect 22657 8002 22658 8036
rect 22802 8010 22803 8021
rect 22646 7968 22647 7979
rect 22813 7976 22814 8010
rect 22969 8002 22970 8036
rect 23114 8010 23115 8021
rect 22958 7968 22959 7979
rect 23125 7976 23126 8010
rect 23281 8002 23282 8036
rect 23270 7968 23271 7979
rect 22345 7934 22346 7968
rect 22490 7942 22491 7953
rect 3082 7908 3083 7919
rect 2135 7874 2136 7908
rect 2447 7874 2448 7908
rect 2759 7874 2760 7908
rect 3071 7874 3072 7908
rect 22334 7900 22335 7911
rect 22501 7908 22502 7942
rect 22657 7934 22658 7968
rect 22802 7942 22803 7953
rect 22646 7900 22647 7911
rect 22813 7908 22814 7942
rect 22969 7934 22970 7968
rect 23114 7942 23115 7953
rect 22958 7900 22959 7911
rect 23125 7908 23126 7942
rect 23281 7934 23282 7968
rect 23270 7900 23271 7911
rect 5036 7870 5051 7898
rect 2146 7702 2147 7713
rect 692 7688 693 7699
rect 1032 7688 1033 7699
rect 1344 7688 1345 7699
rect 1656 7688 1657 7699
rect 681 7654 682 7688
rect 1021 7654 1022 7688
rect 1333 7654 1334 7688
rect 1645 7654 1646 7688
rect 2135 7668 2136 7702
rect 2302 7696 2303 7707
rect 2458 7702 2459 7713
rect 2291 7662 2292 7696
rect 2447 7668 2448 7702
rect 2614 7696 2615 7707
rect 2770 7702 2771 7713
rect 2603 7662 2604 7696
rect 2759 7668 2760 7702
rect 2926 7696 2927 7707
rect 3082 7702 3083 7713
rect 2915 7662 2916 7696
rect 3071 7668 3072 7702
rect 5008 7676 5023 7870
rect 20366 7862 20381 7890
rect 22345 7866 22346 7900
rect 22657 7866 22658 7900
rect 22969 7866 22970 7900
rect 23281 7866 23282 7900
rect 20394 7668 20409 7862
rect 23401 7858 23402 8038
rect 23426 8010 23427 8021
rect 23426 7942 23427 7953
rect 23435 7892 23436 8072
rect 23437 8044 23438 8078
rect 23799 8070 23800 8104
rect 23944 8078 23945 8089
rect 23788 8036 23789 8047
rect 23955 8044 23956 8078
rect 24111 8070 24112 8104
rect 24256 8078 24257 8089
rect 24100 8036 24101 8047
rect 24267 8044 24268 8078
rect 24423 8070 24424 8104
rect 24568 8078 24569 8089
rect 24412 8036 24413 8047
rect 24579 8044 24580 8078
rect 24735 8070 24736 8104
rect 24880 8078 24881 8089
rect 24724 8036 24725 8047
rect 24891 8044 24892 8078
rect 23437 7976 23438 8010
rect 23799 8002 23800 8036
rect 23944 8010 23945 8021
rect 23788 7968 23789 7979
rect 23955 7976 23956 8010
rect 24111 8002 24112 8036
rect 24256 8010 24257 8021
rect 24100 7968 24101 7979
rect 24267 7976 24268 8010
rect 24423 8002 24424 8036
rect 24568 8010 24569 8021
rect 24412 7968 24413 7979
rect 24579 7976 24580 8010
rect 24735 8002 24736 8036
rect 24880 8010 24881 8021
rect 24724 7968 24725 7979
rect 24891 7976 24892 8010
rect 23437 7908 23438 7942
rect 23799 7934 23800 7968
rect 23944 7942 23945 7953
rect 23788 7900 23789 7911
rect 23955 7908 23956 7942
rect 24111 7934 24112 7968
rect 24256 7942 24257 7953
rect 24100 7900 24101 7911
rect 24267 7908 24268 7942
rect 24423 7934 24424 7968
rect 24568 7942 24569 7953
rect 24412 7900 24413 7911
rect 24579 7908 24580 7942
rect 24735 7934 24736 7968
rect 24880 7942 24881 7953
rect 24724 7900 24725 7911
rect 24891 7908 24892 7942
rect 23799 7866 23800 7900
rect 24111 7866 24112 7900
rect 24423 7866 24424 7900
rect 24735 7866 24736 7900
rect 22334 7694 22335 7705
rect 22345 7660 22346 7694
rect 22490 7688 22491 7699
rect 22646 7694 22647 7705
rect 22501 7654 22502 7688
rect 22657 7660 22658 7694
rect 22802 7688 22803 7699
rect 22958 7694 22959 7705
rect 22813 7654 22814 7688
rect 22969 7660 22970 7694
rect 23114 7688 23115 7699
rect 23270 7694 23271 7705
rect 23125 7654 23126 7688
rect 23281 7660 23282 7694
rect 23760 7680 23761 7691
rect 24072 7680 24073 7691
rect 24384 7680 24385 7691
rect 24724 7680 24725 7691
rect 23771 7646 23772 7680
rect 24083 7646 24084 7680
rect 24395 7646 24396 7680
rect 24735 7646 24736 7680
rect 692 7620 693 7631
rect 876 7628 877 7639
rect 681 7586 682 7620
rect 865 7594 866 7628
rect 1032 7620 1033 7631
rect 1188 7628 1189 7639
rect 1021 7586 1022 7620
rect 1177 7594 1178 7628
rect 1344 7620 1345 7631
rect 1500 7628 1501 7639
rect 2146 7634 2147 7645
rect 1333 7586 1334 7620
rect 1489 7594 1490 7628
rect 1656 7620 1657 7631
rect 1645 7586 1646 7620
rect 2135 7600 2136 7634
rect 2302 7628 2303 7639
rect 2458 7634 2459 7645
rect 2291 7594 2292 7628
rect 2447 7600 2448 7634
rect 2614 7628 2615 7639
rect 2770 7634 2771 7645
rect 2603 7594 2604 7628
rect 2759 7600 2760 7634
rect 2926 7628 2927 7639
rect 3082 7634 3083 7645
rect 2915 7594 2916 7628
rect 3071 7600 3072 7634
rect 22334 7626 22335 7637
rect 22345 7592 22346 7626
rect 22490 7620 22491 7631
rect 22646 7626 22647 7637
rect 22501 7586 22502 7620
rect 22657 7592 22658 7626
rect 22802 7620 22803 7631
rect 22958 7626 22959 7637
rect 22813 7586 22814 7620
rect 22969 7592 22970 7626
rect 23114 7620 23115 7631
rect 23270 7626 23271 7637
rect 23125 7586 23126 7620
rect 23281 7592 23282 7626
rect 23760 7612 23761 7623
rect 23916 7620 23917 7631
rect 23771 7578 23772 7612
rect 23927 7586 23928 7620
rect 24072 7612 24073 7623
rect 24228 7620 24229 7631
rect 24083 7578 24084 7612
rect 24239 7586 24240 7620
rect 24384 7612 24385 7623
rect 24540 7620 24541 7631
rect 24395 7578 24396 7612
rect 24551 7586 24552 7620
rect 24724 7612 24725 7623
rect 24735 7578 24736 7612
rect 486 7514 1806 7564
rect 1940 7514 3214 7564
rect 22203 7506 23477 7556
rect 23611 7506 24931 7556
rect 448 7440 3214 7442
rect 22203 7432 24969 7434
rect 894 7132 2498 7182
rect 2510 7132 2710 7182
rect 2796 7132 2996 7182
rect 944 7120 945 7131
rect 1256 7120 1257 7131
rect 1568 7120 1569 7131
rect 1880 7120 1881 7131
rect 2192 7120 2193 7131
rect 2560 7120 2561 7131
rect 933 7086 934 7120
rect 1100 7078 1101 7089
rect 1245 7086 1246 7120
rect 1412 7078 1413 7089
rect 1557 7086 1558 7120
rect 1724 7078 1725 7089
rect 1869 7086 1870 7120
rect 2036 7078 2037 7089
rect 2181 7086 2182 7120
rect 2348 7078 2349 7089
rect 2549 7086 2550 7120
rect 2945 7086 2946 7131
rect 22421 7124 22621 7174
rect 22707 7124 22907 7174
rect 22919 7124 24523 7174
rect 22471 7078 22472 7123
rect 22856 7112 22857 7123
rect 23224 7112 23225 7123
rect 23536 7112 23537 7123
rect 23848 7112 23849 7123
rect 24160 7112 24161 7123
rect 24472 7112 24473 7123
rect 22867 7078 22868 7112
rect 944 7052 945 7063
rect 933 7018 934 7052
rect 1089 7044 1090 7078
rect 1256 7052 1257 7063
rect 1100 7010 1101 7021
rect 1245 7018 1246 7052
rect 1401 7044 1402 7078
rect 1568 7052 1569 7063
rect 1412 7010 1413 7021
rect 1557 7018 1558 7052
rect 1713 7044 1714 7078
rect 1880 7052 1881 7063
rect 1724 7010 1725 7021
rect 1869 7018 1870 7052
rect 2025 7044 2026 7078
rect 2192 7052 2193 7063
rect 2036 7010 2037 7021
rect 2181 7018 2182 7052
rect 2337 7044 2338 7078
rect 23068 7070 23069 7081
rect 23235 7078 23236 7112
rect 23380 7070 23381 7081
rect 23547 7078 23548 7112
rect 23692 7070 23693 7081
rect 23859 7078 23860 7112
rect 24004 7070 24005 7081
rect 24171 7078 24172 7112
rect 24316 7070 24317 7081
rect 24483 7078 24484 7112
rect 2560 7052 2561 7063
rect 2348 7010 2349 7021
rect 2549 7018 2550 7052
rect 2945 7012 2946 7057
rect 944 6984 945 6995
rect 933 6950 934 6984
rect 1089 6976 1090 7010
rect 1256 6984 1257 6995
rect 1100 6942 1101 6953
rect 1245 6950 1246 6984
rect 1401 6976 1402 7010
rect 1568 6984 1569 6995
rect 1412 6942 1413 6953
rect 1557 6950 1558 6984
rect 1713 6976 1714 7010
rect 1880 6984 1881 6995
rect 1724 6942 1725 6953
rect 1869 6950 1870 6984
rect 2025 6976 2026 7010
rect 2192 6984 2193 6995
rect 2036 6942 2037 6953
rect 2181 6950 2182 6984
rect 2337 6976 2338 7010
rect 3116 7002 3214 7052
rect 2560 6984 2561 6995
rect 22203 6994 22301 7044
rect 22471 7004 22472 7049
rect 22856 7044 22857 7055
rect 22867 7010 22868 7044
rect 23079 7036 23080 7070
rect 23224 7044 23225 7055
rect 23068 7002 23069 7013
rect 23235 7010 23236 7044
rect 23391 7036 23392 7070
rect 23536 7044 23537 7055
rect 23380 7002 23381 7013
rect 23547 7010 23548 7044
rect 23703 7036 23704 7070
rect 23848 7044 23849 7055
rect 23692 7002 23693 7013
rect 23859 7010 23860 7044
rect 24015 7036 24016 7070
rect 24160 7044 24161 7055
rect 24004 7002 24005 7013
rect 24171 7010 24172 7044
rect 24327 7036 24328 7070
rect 24472 7044 24473 7055
rect 24316 7002 24317 7013
rect 24483 7010 24484 7044
rect 2348 6942 2349 6953
rect 2549 6950 2550 6984
rect 944 6916 945 6927
rect 933 6882 934 6916
rect 935 6866 936 6916
rect 1089 6908 1090 6942
rect 1256 6916 1257 6927
rect 969 6832 970 6882
rect 1100 6874 1101 6885
rect 1245 6882 1246 6916
rect 1401 6908 1402 6942
rect 1568 6916 1569 6927
rect 1412 6874 1413 6885
rect 1557 6882 1558 6916
rect 1713 6908 1714 6942
rect 1880 6916 1881 6927
rect 1724 6874 1725 6885
rect 1869 6882 1870 6916
rect 2025 6908 2026 6942
rect 2192 6916 2193 6927
rect 2036 6874 2037 6885
rect 2181 6882 2182 6916
rect 2337 6908 2338 6942
rect 2945 6938 2946 6983
rect 22856 6976 22857 6987
rect 22471 6930 22472 6975
rect 22867 6942 22868 6976
rect 23079 6968 23080 7002
rect 23224 6976 23225 6987
rect 23068 6934 23069 6945
rect 23235 6942 23236 6976
rect 23391 6968 23392 7002
rect 23536 6976 23537 6987
rect 23380 6934 23381 6945
rect 23547 6942 23548 6976
rect 23703 6968 23704 7002
rect 23848 6976 23849 6987
rect 23692 6934 23693 6945
rect 23859 6942 23860 6976
rect 24015 6968 24016 7002
rect 24160 6976 24161 6987
rect 24004 6934 24005 6945
rect 24171 6942 24172 6976
rect 24327 6968 24328 7002
rect 24472 6976 24473 6987
rect 24316 6934 24317 6945
rect 24483 6942 24484 6976
rect 2560 6916 2561 6927
rect 2348 6874 2349 6885
rect 2549 6882 2550 6916
rect 22856 6908 22857 6919
rect 1089 6840 1090 6874
rect 1401 6840 1402 6874
rect 1713 6840 1714 6874
rect 2025 6840 2026 6874
rect 2337 6840 2338 6874
rect 2945 6860 2946 6905
rect 22471 6852 22472 6897
rect 22867 6874 22868 6908
rect 23079 6900 23080 6934
rect 23224 6908 23225 6919
rect 23068 6866 23069 6877
rect 23235 6874 23236 6908
rect 23391 6900 23392 6934
rect 23536 6908 23537 6919
rect 23380 6866 23381 6877
rect 23547 6874 23548 6908
rect 23703 6900 23704 6934
rect 23848 6908 23849 6919
rect 23692 6866 23693 6877
rect 23859 6874 23860 6908
rect 24015 6900 24016 6934
rect 24160 6908 24161 6919
rect 24004 6866 24005 6877
rect 24171 6874 24172 6908
rect 24327 6900 24328 6934
rect 24472 6908 24473 6919
rect 24316 6866 24317 6877
rect 3116 6802 3214 6852
rect 22203 6794 22301 6844
rect 23079 6832 23080 6866
rect 23391 6832 23392 6866
rect 23703 6832 23704 6866
rect 24015 6832 24016 6866
rect 24327 6832 24328 6866
rect 24447 6824 24448 6874
rect 24481 6858 24482 6908
rect 24483 6874 24484 6908
rect 1100 6668 1101 6679
rect 1089 6634 1090 6668
rect 1256 6662 1257 6673
rect 1412 6668 1413 6679
rect 1245 6628 1246 6662
rect 1401 6634 1402 6668
rect 1568 6662 1569 6673
rect 1724 6668 1725 6679
rect 1557 6628 1558 6662
rect 1713 6634 1714 6668
rect 1880 6662 1881 6673
rect 2036 6668 2037 6679
rect 1869 6628 1870 6662
rect 2025 6634 2026 6668
rect 2192 6662 2193 6673
rect 2181 6628 2182 6662
rect 2348 6654 2349 6665
rect 2337 6620 2338 6654
rect 23068 6646 23069 6657
rect 23224 6654 23225 6665
rect 23380 6660 23381 6671
rect 1100 6600 1101 6611
rect 1089 6566 1090 6600
rect 1256 6594 1257 6605
rect 1412 6600 1413 6611
rect 1245 6560 1246 6594
rect 1401 6566 1402 6600
rect 1568 6594 1569 6605
rect 1724 6600 1725 6611
rect 1557 6560 1558 6594
rect 1713 6566 1714 6600
rect 1880 6594 1881 6605
rect 2036 6600 2037 6611
rect 1869 6560 1870 6594
rect 2025 6566 2026 6600
rect 2192 6594 2193 6605
rect 2181 6560 2182 6594
rect 2348 6586 2349 6597
rect 2945 6596 2946 6641
rect 2337 6552 2338 6586
rect 894 6480 2498 6530
rect 2506 6480 2706 6530
rect 2945 6528 2946 6573
rect 3162 6564 3214 6614
rect 22203 6556 22255 6606
rect 22471 6588 22472 6633
rect 23079 6612 23080 6646
rect 23235 6620 23236 6654
rect 23391 6626 23392 6660
rect 23536 6654 23537 6665
rect 23692 6660 23693 6671
rect 23547 6620 23548 6654
rect 23703 6626 23704 6660
rect 23848 6654 23849 6665
rect 24004 6660 24005 6671
rect 23859 6620 23860 6654
rect 24015 6626 24016 6660
rect 24160 6654 24161 6665
rect 24316 6660 24317 6671
rect 24171 6620 24172 6654
rect 24327 6626 24328 6660
rect 23068 6578 23069 6589
rect 23224 6586 23225 6597
rect 23380 6592 23381 6603
rect 22471 6520 22472 6565
rect 23079 6544 23080 6578
rect 23235 6552 23236 6586
rect 23391 6558 23392 6592
rect 23536 6586 23537 6597
rect 23692 6592 23693 6603
rect 23547 6552 23548 6586
rect 23703 6558 23704 6592
rect 23848 6586 23849 6597
rect 24004 6592 24005 6603
rect 23859 6552 23860 6586
rect 24015 6558 24016 6592
rect 24160 6586 24161 6597
rect 24316 6592 24317 6603
rect 24171 6552 24172 6586
rect 24327 6558 24328 6592
rect 2796 6446 2996 6496
rect 22421 6438 22621 6488
rect 22711 6472 22911 6522
rect 22919 6472 24523 6522
rect 490 6406 524 6408
rect 586 6406 620 6408
rect 682 6406 716 6408
rect 778 6406 812 6408
rect 874 6406 908 6408
rect 970 6406 1004 6408
rect 1066 6406 1100 6408
rect 1162 6406 1196 6408
rect 1258 6406 1292 6408
rect 1354 6406 1388 6408
rect 1450 6406 1484 6408
rect 1546 6406 1580 6408
rect 1642 6406 1676 6408
rect 1738 6406 1772 6408
rect 1834 6406 1868 6408
rect 1930 6406 1964 6408
rect 2026 6406 2060 6408
rect 2122 6406 2156 6408
rect 2218 6406 2252 6408
rect 2314 6406 2348 6408
rect 2410 6406 2444 6408
rect 2506 6406 2540 6408
rect 2602 6406 2636 6408
rect 2698 6406 2732 6408
rect 2794 6406 2828 6408
rect 2890 6406 2924 6408
rect 2986 6406 3020 6408
rect 3082 6406 3116 6408
rect 3178 6406 3212 6408
rect 22205 6398 22239 6400
rect 22301 6398 22335 6400
rect 22397 6398 22431 6400
rect 22493 6398 22527 6400
rect 22589 6398 22623 6400
rect 22685 6398 22719 6400
rect 22781 6398 22815 6400
rect 22877 6398 22911 6400
rect 22973 6398 23007 6400
rect 23069 6398 23103 6400
rect 23165 6398 23199 6400
rect 23261 6398 23295 6400
rect 23357 6398 23391 6400
rect 23453 6398 23487 6400
rect 23549 6398 23583 6400
rect 23645 6398 23679 6400
rect 23741 6398 23775 6400
rect 23837 6398 23871 6400
rect 23933 6398 23967 6400
rect 24029 6398 24063 6400
rect 24125 6398 24159 6400
rect 24221 6398 24255 6400
rect 24317 6398 24351 6400
rect 24413 6398 24447 6400
rect 24509 6398 24543 6400
rect 24605 6398 24639 6400
rect 24701 6398 24735 6400
rect 24797 6398 24831 6400
rect 24893 6398 24927 6400
use example_por  example_por_0
timestamp 1695321174
transform -1 0 11285 0 1 -14
box 0 0 11344 8338
use example_por  example_por_1
timestamp 1695321174
transform 1 0 14132 0 1 -22
box 0 0 11344 8338
<< end >>

* NGSPICE file created from ldo.ext - technology: sky130A

.subckt ldo Iref VB VS OUT SS DD
X0 a_9110_n8196.t3 VB.t0 a_8766_n8196.t1 SS.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=5.19 l=1.43
X1 SS.t1 Iref.t4 a_9110_n8196.t0 SS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X2 DD.t7 a_8766_n8196.t4 OUT.t3 DD.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.9 as=1.5 ps=10.9 w=5.17 l=0.37
X3 DD.t15 DD.t12 DD.t14 DD.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.258 ps=2.36 w=0.89 l=3.89
X4 a_9110_n8196.t6 Iref.t5 SS.t22 SS.t21 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X5 a_8766_n8196.t5 OUT.t2 sky130_fd_pr__cap_mim_m3_1 l=15 w=4
X6 DD.t17 a_9330_n9998.t4 a_9330_n9998.t5 DD.t16 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X7 DD.t5 a_9330_n9998.t6 a_8766_n8196.t3 DD.t4 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X8 SS.t6 Iref.t6 a_9330_n9998.t1 SS.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X9 SS.t20 SS.t17 SS.t19 SS.t18 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=1.48 ps=10.8 w=5.1 l=0.66
X10 OUT.t4 VS.t0 a_9110_n8196.t7 OUT.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.76 pd=12.7 as=1.76 ps=12.7 w=6.07 l=1.27
X11 a_9110_n8196.t4 Iref.t7 SS.t8 SS.t7 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X12 SS.t24 Iref.t2 Iref.t3 SS.t23 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X13 DD.t1 a_9330_n9998.t7 a_8766_n8196.t0 DD.t0 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X14 OUT.t1 VS.t1 a_9110_n8196.t1 OUT.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.76 pd=12.7 as=1.76 ps=12.7 w=6.07 l=1.27
X15 SS.t12 Iref.t8 a_9110_n8196.t5 SS.t11 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X16 a_9110_n8196.t2 VB.t1 a_8766_n8196.t2 SS.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.51 pd=11 as=1.51 ps=11 w=5.19 l=1.43
X17 DD.t11 DD.t8 DD.t10 DD.t9 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0 ps=0 w=0.89 l=3.89
X18 SS.t16 SS.t13 SS.t15 SS.t14 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=0 ps=0 w=5.1 l=0.66
X19 DD.t3 a_9330_n9998.t2 a_9330_n9998.t3 DD.t2 sky130_fd_pr__pfet_01v8 ad=0.258 pd=2.36 as=0.258 ps=2.36 w=0.89 l=3.89
X20 a_9330_n9998.t0 Iref.t9 SS.t3 SS.t2 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
X21 Iref.t1 Iref.t0 SS.t10 SS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.48 pd=10.8 as=1.48 ps=10.8 w=5.1 l=0.66
R0 VB.n0 VB.t0 49.9518
R1 VB.n0 VB.t1 48.1905
R2 VB VB.n0 2.76135
R3 a_8766_n8196.n0 a_8766_n8196.t4 191.636
R4 a_8766_n8196.n0 a_8766_n8196.t0 34.661
R5 a_8766_n8196.n0 a_8766_n8196.t3 33.291
R6 a_8766_n8196.t1 a_8766_n8196.n1 4.51459
R7 a_8766_n8196.n1 a_8766_n8196.t2 3.35375
R8 a_8766_n8196.t5 a_8766_n8196.n0 2.51069
R9 a_8766_n8196.n1 a_8766_n8196.t5 1.37236
R10 a_9110_n8196.n0 a_9110_n8196.t7 7.40825
R11 a_9110_n8196.n0 a_9110_n8196.t1 4.70699
R12 a_9110_n8196.n1 a_9110_n8196.t5 4.53569
R13 a_9110_n8196.n3 a_9110_n8196.t4 4.53369
R14 a_9110_n8196.n4 a_9110_n8196.t6 4.38957
R15 a_9110_n8196.t0 a_9110_n8196.n5 4.3873
R16 a_9110_n8196.n2 a_9110_n8196.t2 4.26166
R17 a_9110_n8196.n2 a_9110_n8196.t3 4.06962
R18 a_9110_n8196.n5 a_9110_n8196.n4 2.26478
R19 a_9110_n8196.n3 a_9110_n8196.n2 2.0915
R20 a_9110_n8196.n1 a_9110_n8196.n0 0.66715
R21 a_9110_n8196.n4 a_9110_n8196.n3 0.1505
R22 a_9110_n8196.n5 a_9110_n8196.n1 0.144506
R23 SS.n18 SS.n17 4862.2
R24 SS.n8 SS.n6 1303.68
R25 SS.t14 SS.t5 969.697
R26 SS.t0 SS.t11 969.697
R27 SS.n20 SS.n16 774.62
R28 SS.n9 SS.n1 770.619
R29 SS.n23 SS.t14 623.03
R30 SS.n1 SS.n0 610.112
R31 SS.n24 SS.n22 604.529
R32 SS.n28 SS.t0 438.788
R33 SS.n16 SS.n13 380.226
R34 SS.t9 SS.t21 344.896
R35 SS.t2 SS.t7 344.896
R36 SS.n19 SS.n18 293.863
R37 SS.n26 SS.n20 280.995
R38 SS.n40 SS.n27 270.781
R39 SS.t4 SS.n4 246.601
R40 SS.n41 SS.n40 227.38
R41 SS.n11 SS.t16 220.899
R42 SS.n29 SS.t13 220.834
R43 SS.n42 SS.t19 220.522
R44 SS.n42 SS.t17 206.317
R45 SS.n38 SS.t9 193.142
R46 SS.t23 SS.n28 188.831
R47 SS.n38 SS.t23 151.755
R48 SS.n30 SS.t6 127.653
R49 SS.n31 SS.t12 127.653
R50 SS.n32 SS.t1 127.653
R51 SS.n33 SS.t24 127.653
R52 SS.n35 SS.t10 127.653
R53 SS.n34 SS.t22 127.653
R54 SS.n47 SS.t8 127.653
R55 SS.n48 SS.t3 127.653
R56 SS.n50 SS.n49 119.424
R57 SS.n52 SS.n51 102.663
R58 SS.t4 SS.t18 88.811
R59 SS.n27 SS.n26 72.8795
R60 SS.t18 SS.n5 64.6683
R61 SS.n31 SS.n30 60.9529
R62 SS.n32 SS.n31 60.9529
R63 SS.n33 SS.n32 60.9529
R64 SS.n35 SS.n34 60.9529
R65 SS.n48 SS.n47 60.9529
R66 SS.n46 SS.n45 56.9082
R67 SS.n36 SS.n35 54.7053
R68 SS.n36 SS.n33 47.2386
R69 SS.n30 SS.n29 40.3815
R70 SS.n49 SS.n48 40.0767
R71 SS.n26 SS.n25 22.3606
R72 SS.n27 SS.n11 17.6395
R73 SS.n52 SS.n42 17.6395
R74 SS.n4 SS.t2 9.48512
R75 SS.n21 SS.t15 3.47896
R76 SS.n50 SS.t20 3.41269
R77 SS SS.n41 2.09505
R78 SS.n41 SS.n10 1.88285
R79 SS.n51 SS.n50 1.38918
R80 SS SS.n52 0.756864
R81 SS.n25 SS.n21 0.126275
R82 SS.n25 SS.n24 0.100882
R83 SS.n10 SS.n9 0.0360926
R84 SS.n9 SS.t4 0.0360926
R85 SS.n8 SS.n7 0.0360926
R86 SS.t4 SS.n8 0.0360926
R87 SS.n3 SS.n2 0.00609809
R88 SS.n4 SS.n3 0.00609809
R89 SS.n44 SS.n43 0.00609809
R90 SS.n45 SS.n44 0.00609809
R91 SS.n16 SS.n15 0.00100268
R92 SS.n24 SS.n23 0.00051152
R93 SS.n51 SS.n46 0.00051152
R94 SS.n13 SS.n12 0.000510263
R95 SS.n40 SS.n39 0.000503106
R96 SS.n39 SS.n38 0.000503106
R97 SS.n38 SS.n37 0.000503106
R98 SS.n37 SS.n36 0.000503106
R99 SS.n15 SS.n14 0.000502681
R100 SS.n20 SS.n19 0.000501887
R101 Iref.n10 Iref.t9 206.963
R102 Iref.n2 Iref.t6 206.963
R103 Iref.n2 Iref.t8 206.321
R104 Iref.n4 Iref.t4 206.321
R105 Iref.n6 Iref.t2 206.321
R106 Iref.n10 Iref.t7 206.321
R107 Iref.n11 Iref.t5 206.321
R108 Iref.n12 Iref.t0 206.321
R109 Iref.t8 Iref.n1 206.317
R110 Iref.t4 Iref.n3 206.317
R111 Iref.t2 Iref.n5 206.317
R112 Iref.t7 Iref.n9 206.317
R113 Iref.t5 Iref.n8 206.317
R114 Iref.t0 Iref.n7 206.317
R115 Iref.n0 Iref.t1 3.41293
R116 Iref.n0 Iref.t3 3.41293
R117 Iref.n12 Iref.n11 0.642396
R118 Iref.n11 Iref.n10 0.642396
R119 Iref.n4 Iref.n2 0.642396
R120 Iref.n6 Iref.n4 0.642396
R121 Iref.n13 Iref.n12 0.237335
R122 Iref.n13 Iref.n6 0.235494
R123 Iref Iref.n13 0.20576
R124 Iref Iref.n0 0.184094
R125 OUT.n9 OUT.n8 261.185
R126 OUT.n4 OUT.n3 229.173
R127 OUT.n12 OUT.n11 74.0415
R128 OUT.n12 OUT.n6 72.1843
R129 OUT.n1 OUT.t1 7.2144
R130 OUT.n25 OUT.t3 5.76538
R131 OUT.n0 OUT.t4 4.7068
R132 OUT.n19 OUT.t0 4.24157
R133 OUT.n13 OUT.n12 1.23559
R134 OUT OUT.n25 0.180481
R135 OUT.n24 OUT.n23 0.136226
R136 OUT.n24 OUT.t2 0.126657
R137 OUT.n14 OUT.n1 0.0503555
R138 OUT.n23 OUT.n14 0.0427877
R139 OUT.n1 OUT.n0 0.0245405
R140 OUT.n25 OUT.n24 0.0179077
R141 OUT.n6 OUT.n5 0.0153511
R142 OUT.n5 OUT.n4 0.014836
R143 OUT.n11 OUT.n10 0.0131168
R144 OUT.n10 OUT.n9 0.012684
R145 OUT.n21 OUT.n20 0.0069195
R146 OUT.n20 OUT.n19 0.00641981
R147 OUT.n23 OUT.n22 0.00626716
R148 OUT.n21 OUT.n16 0.00449474
R149 OUT.n8 OUT.n7 0.00432563
R150 OUT.n3 OUT.n2 0.00432563
R151 OUT.n16 OUT.n15 0.00399493
R152 OUT.n18 OUT.n17 0.00345991
R153 OUT.n19 OUT.n18 0.00345991
R154 OUT.n22 OUT.n21 0.00100012
R155 OUT.n14 OUT.n13 0.000504061
R156 DD.n3 DD.n2 459.671
R157 DD.t9 DD.t4 367.363
R158 DD.t16 DD.t0 367.363
R159 DD.n26 DD.n20 282.247
R160 DD.n9 DD.n8 254.948
R161 DD.n0 DD.t9 232.912
R162 DD.n7 DD.t13 213.075
R163 DD.n27 DD.n18 209.695
R164 DD.n5 DD.t16 193.233
R165 DD.n16 DD.n15 186.632
R166 DD.n5 DD.t2 174.131
R167 DD.n29 DD.n27 63.0245
R168 DD.n2 DD.t15 60.0995
R169 DD.n28 DD.t11 60.0995
R170 DD.n29 DD.n28 53.4946
R171 DD.n9 DD.t14 48.3828
R172 DD.n15 DD.t10 45.276
R173 DD.n14 DD.n13 34.174
R174 DD.n11 DD.n10 34.174
R175 DD.n10 DD.t1 32.0995
R176 DD.n11 DD.t17 32.0995
R177 DD.n13 DD.t3 32.0995
R178 DD.n14 DD.t5 32.0995
R179 DD.n15 DD.n14 28.5054
R180 DD.n10 DD.n9 28.5054
R181 DD.n12 DD.n11 18.0327
R182 DD.n13 DD.n12 16.1418
R183 DD.n27 DD.n26 10.8113
R184 DD.n1 DD.t8 9.47999
R185 DD.n8 DD.t12 9.47999
R186 DD.n30 DD.n29 8.40959
R187 DD.n31 DD.n16 8.10924
R188 DD.n26 DD.t7 5.52608
R189 DD.n31 DD.n30 5.40633
R190 DD.n16 DD.n1 0.840904
R191 DD DD.n31 0.196382
R192 DD.n18 DD.n17 0.025954
R193 DD.n20 DD.n19 0.025954
R194 DD.n8 DD.n7 0.00450849
R195 DD.n1 DD.n0 0.00450849
R196 DD.n22 DD.n21 0.00414317
R197 DD.n26 DD.n25 0.00414317
R198 DD.n25 DD.n24 0.00355895
R199 DD.n23 DD.n22 0.00348454
R200 DD.n24 DD.t6 0.00231816
R201 DD.t6 DD.n23 0.00215862
R202 DD.n12 DD.n6 0.00193193
R203 DD.n6 DD.n5 0.00193193
R204 DD.n5 DD.n4 0.00193193
R205 DD.n4 DD.n3 0.00193193
R206 a_9330_n9998.n1 a_9330_n9998.t5 32.4466
R207 a_9330_n9998.n0 a_9330_n9998.t3 32.4466
R208 a_9330_n9998.t4 a_9330_n9998.t7 19.1411
R209 a_9330_n9998.t2 a_9330_n9998.t6 19.1411
R210 a_9330_n9998.t1 a_9330_n9998.n4 10.1828
R211 a_9330_n9998.n3 a_9330_n9998.t4 9.48031
R212 a_9330_n9998.n2 a_9330_n9998.t2 9.48031
R213 a_9330_n9998.n4 a_9330_n9998.n1 5.92365
R214 a_9330_n9998.n4 a_9330_n9998.t0 5.36911
R215 a_9330_n9998.n0 a_9330_n9998.n2 0.351043
R216 a_9330_n9998.n1 a_9330_n9998.n3 0.351043
R217 a_9330_n9998.n1 a_9330_n9998.n0 0.100294
R218 VS.n0 VS.t1 147.147
R219 VS.n0 VS.t0 63.6678
R220 VS VS.n0 44.4531
C0 Iref VB 0.267f
C1 OUT DD 1.36f
C2 DD VS 0.00151f
C3 OUT VS 2.33f
C4 OUT Iref 0.0248f
C5 DD VB 0.0106f
C6 Iref VS 0.00227f
C7 OUT VB 1.46f
C8 VB VS 0.134f
.ends


magic
tech sky130A
timestamp 1695672277
<< nmoslvt >>
rect -50 -275 50 275
<< ndiff >>
rect -79 269 -50 275
rect -79 -269 -73 269
rect -56 -269 -50 269
rect -79 -275 -50 -269
rect 50 269 79 275
rect 50 -269 56 269
rect 73 -269 79 269
rect 50 -275 79 -269
<< ndiffc >>
rect -73 -269 -56 269
rect 56 -269 73 269
<< poly >>
rect -50 311 50 319
rect -50 294 -42 311
rect 42 294 50 311
rect -50 275 50 294
rect -50 -294 50 -275
rect -50 -311 -42 -294
rect 42 -311 50 -294
rect -50 -319 50 -311
<< polycont >>
rect -42 294 42 311
rect -42 -311 42 -294
<< locali >>
rect -50 294 -42 311
rect 42 294 50 311
rect -73 269 -56 277
rect -73 -277 -56 -269
rect 56 269 73 277
rect 56 -277 73 -269
rect -50 -311 -42 -294
rect 42 -311 50 -294
<< viali >>
rect -42 294 42 311
rect -73 -269 -56 269
rect 56 -269 73 269
rect -42 -311 42 -294
<< metal1 >>
rect -48 311 48 314
rect -48 294 -42 311
rect 42 294 48 311
rect -48 291 48 294
rect -76 269 -53 275
rect -76 -269 -73 269
rect -56 -269 -53 269
rect -76 -275 -53 -269
rect 53 269 76 275
rect 53 -269 56 269
rect 73 -269 76 269
rect 53 -275 76 -269
rect -48 -294 48 -291
rect -48 -311 -42 -294
rect 42 -311 48 -294
rect -48 -314 48 -311
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.5 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

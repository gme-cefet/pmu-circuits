magic
tech sky130A
magscale 1 2
timestamp 1696345916
<< pwell >>
rect -339 -1357 339 1357
<< nmoslvt >>
rect -143 109 143 1147
rect -143 -1147 143 -109
<< ndiff >>
rect -201 1135 -143 1147
rect -201 121 -189 1135
rect -155 121 -143 1135
rect -201 109 -143 121
rect 143 1135 201 1147
rect 143 121 155 1135
rect 189 121 201 1135
rect 143 109 201 121
rect -201 -121 -143 -109
rect -201 -1135 -189 -121
rect -155 -1135 -143 -121
rect -201 -1147 -143 -1135
rect 143 -121 201 -109
rect 143 -1135 155 -121
rect 189 -1135 201 -121
rect 143 -1147 201 -1135
<< ndiffc >>
rect -189 121 -155 1135
rect 155 121 189 1135
rect -189 -1135 -155 -121
rect 155 -1135 189 -121
<< psubdiff >>
rect -303 1287 -207 1321
rect 207 1287 303 1321
rect -303 1225 -269 1287
rect 269 1225 303 1287
rect -303 -1287 -269 -1225
rect 269 -1287 303 -1225
rect -303 -1321 -207 -1287
rect 207 -1321 303 -1287
<< psubdiffcont >>
rect -207 1287 207 1321
rect -303 -1225 -269 1225
rect 269 -1225 303 1225
rect -207 -1321 207 -1287
<< poly >>
rect -143 1219 143 1235
rect -143 1185 -127 1219
rect 127 1185 143 1219
rect -143 1147 143 1185
rect -143 71 143 109
rect -143 37 -127 71
rect 127 37 143 71
rect -143 21 143 37
rect -143 -37 143 -21
rect -143 -71 -127 -37
rect 127 -71 143 -37
rect -143 -109 143 -71
rect -143 -1185 143 -1147
rect -143 -1219 -127 -1185
rect 127 -1219 143 -1185
rect -143 -1235 143 -1219
<< polycont >>
rect -127 1185 127 1219
rect -127 37 127 71
rect -127 -71 127 -37
rect -127 -1219 127 -1185
<< locali >>
rect -303 1287 -207 1321
rect 207 1287 303 1321
rect -303 1225 -269 1287
rect 269 1225 303 1287
rect -143 1185 -127 1219
rect 127 1185 143 1219
rect -189 1135 -155 1151
rect -189 105 -155 121
rect 155 1135 189 1151
rect 155 105 189 121
rect -143 37 -127 71
rect 127 37 143 71
rect -143 -71 -127 -37
rect 127 -71 143 -37
rect -189 -121 -155 -105
rect -189 -1151 -155 -1135
rect 155 -121 189 -105
rect 155 -1151 189 -1135
rect -143 -1219 -127 -1185
rect 127 -1219 143 -1185
rect -303 -1287 -269 -1225
rect 269 -1287 303 -1225
rect -303 -1321 -207 -1287
rect 207 -1321 303 -1287
<< viali >>
rect -127 1185 127 1219
rect -189 121 -155 1135
rect 155 121 189 1135
rect -127 37 127 71
rect -127 -71 127 -37
rect -189 -1135 -155 -121
rect 155 -1135 189 -121
rect -127 -1219 127 -1185
<< metal1 >>
rect -139 1219 139 1225
rect -139 1185 -127 1219
rect 127 1185 139 1219
rect -139 1179 139 1185
rect -195 1135 -149 1147
rect -195 121 -189 1135
rect -155 121 -149 1135
rect -195 109 -149 121
rect 149 1135 195 1147
rect 149 121 155 1135
rect 189 121 195 1135
rect 149 109 195 121
rect -139 71 139 77
rect -139 37 -127 71
rect 127 37 139 71
rect -139 31 139 37
rect -139 -37 139 -31
rect -139 -71 -127 -37
rect 127 -71 139 -37
rect -139 -77 139 -71
rect -195 -121 -149 -109
rect -195 -1135 -189 -121
rect -155 -1135 -149 -121
rect -195 -1147 -149 -1135
rect 149 -121 195 -109
rect 149 -1135 155 -121
rect 189 -1135 195 -121
rect 149 -1147 195 -1135
rect -139 -1185 139 -1179
rect -139 -1219 -127 -1185
rect 127 -1219 139 -1185
rect -139 -1225 139 -1219
<< properties >>
string FIXED_BBOX -286 -1304 286 1304
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.19 l 1.43 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

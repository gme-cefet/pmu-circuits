magic
tech sky130A
magscale 1 2
timestamp 1697038384
<< nwell >>
rect 6759 -3211 10089 -2213
<< psubdiff >>
rect 3175 -164 3305 -140
rect 10257 -164 10387 -140
rect 3305 -315 3377 -191
rect 10166 -315 10257 -191
rect 3305 -3738 3370 -3614
rect 10159 -3738 10257 -3614
rect 3175 -3762 3305 -3738
rect 10257 -3762 10387 -3738
<< nsubdiff >>
rect 6823 -2295 6883 -2261
rect 7937 -2295 7997 -2261
rect 6823 -2321 6857 -2295
rect 6823 -3043 6857 -3017
rect 7963 -2321 7997 -2295
rect 7963 -3043 7997 -3017
rect 6823 -3077 6883 -3043
rect 7937 -3077 7997 -3043
rect 8116 -2306 8176 -2272
rect 9959 -2306 10019 -2272
rect 8116 -2332 8150 -2306
rect 8116 -3123 8150 -3097
rect 9985 -2332 10019 -2306
rect 9985 -3123 10019 -3097
rect 8116 -3157 8176 -3123
rect 9959 -3157 10019 -3123
<< psubdiffcont >>
rect 3175 -3738 3305 -164
rect 3377 -315 10166 -191
rect 3370 -3738 10159 -3614
rect 10257 -3738 10387 -164
<< nsubdiffcont >>
rect 6883 -2295 7937 -2261
rect 6823 -3017 6857 -2321
rect 7963 -3017 7997 -2321
rect 6883 -3077 7937 -3043
rect 8176 -2306 9959 -2272
rect 8116 -3097 8150 -2332
rect 9985 -3097 10019 -2332
rect 8176 -3157 9959 -3123
<< locali >>
rect 3175 -164 3305 -148
rect 10257 -164 10387 -148
rect 3305 -315 3377 -191
rect 10166 -315 10257 -191
rect 4700 -372 4828 -315
rect 8004 -372 8096 -315
rect 4700 -396 8096 -372
rect 3392 -541 3910 -506
rect 3392 -544 9766 -541
rect 3392 -1777 3444 -544
rect 3606 -575 9766 -544
rect 3606 -1777 9766 -1751
rect 3392 -1785 9766 -1777
rect 3392 -1815 3908 -1785
rect 7789 -2034 7962 -1785
rect 7784 -2065 8276 -2034
rect 7784 -2162 7825 -2065
rect 8240 -2162 8276 -2065
rect 7784 -2182 8276 -2162
rect 6626 -2204 6678 -2203
rect 3485 -2252 6678 -2204
rect 3485 -2275 6393 -2252
rect 3485 -3470 6429 -3451
rect 6626 -3470 6678 -2252
rect 6823 -2295 6883 -2261
rect 7937 -2278 7997 -2261
rect 8116 -2278 8176 -2272
rect 7937 -2295 8176 -2278
rect 6823 -2321 6857 -2295
rect 7963 -2306 8176 -2295
rect 9959 -2306 10019 -2272
rect 7963 -2321 8150 -2306
rect 6957 -2462 7252 -2461
rect 6944 -2503 7252 -2462
rect 6944 -2820 6989 -2503
rect 7289 -2519 7529 -2485
rect 7316 -2768 7501 -2718
rect 6944 -2862 7266 -2820
rect 6944 -2864 6989 -2862
rect 6823 -3043 6857 -3017
rect 7384 -3043 7436 -2768
rect 7997 -2332 8150 -2321
rect 7997 -3017 8116 -2332
rect 7963 -3043 8116 -3017
rect 6823 -3077 6883 -3043
rect 7937 -3056 8116 -3043
rect 7937 -3077 7997 -3056
rect 9985 -2332 10019 -2306
rect 8388 -2548 9748 -2514
rect 8644 -2842 8692 -2548
rect 9440 -2842 9488 -2548
rect 8388 -2876 9748 -2842
rect 8116 -3123 8150 -3097
rect 8865 -3029 9258 -3013
rect 8865 -3118 8895 -3029
rect 9235 -3118 9258 -3029
rect 8865 -3123 9258 -3118
rect 9985 -3123 10019 -3097
rect 8116 -3157 8176 -3123
rect 9959 -3157 10019 -3123
rect 8224 -3188 8526 -3157
rect 6725 -3407 7342 -3375
rect 6725 -3470 6767 -3407
rect 3485 -3505 6767 -3470
rect 7309 -3505 7342 -3407
rect 3485 -3525 7342 -3505
rect 6725 -3537 7342 -3525
rect 8224 -3503 8261 -3188
rect 8486 -3503 8526 -3188
rect 8224 -3540 8526 -3503
rect 4134 -3614 5736 -3587
rect 3305 -3738 3370 -3614
rect 10159 -3738 10257 -3614
rect 3175 -3754 3305 -3738
rect 10257 -3754 10387 -3738
<< viali >>
rect 4828 -315 8004 -236
rect 4828 -372 8004 -315
rect 7825 -2162 8240 -2065
rect 8895 -3118 9235 -3029
rect 6767 -3505 7309 -3407
rect 8261 -3503 8486 -3188
rect 4192 -3715 5698 -3616
<< metal1 >>
rect 4700 -236 8096 -200
rect 4700 -372 4828 -236
rect 8004 -372 8096 -236
rect 4700 -377 8096 -372
rect 3512 -410 9554 -377
rect 3512 -1713 3554 -410
rect 3818 -1885 3860 -613
rect 3912 -1713 3954 -410
rect 4218 -1885 4260 -613
rect 4312 -1713 4354 -410
rect 4618 -1885 4660 -613
rect 4712 -1713 4754 -410
rect 5018 -1885 5060 -613
rect 5112 -1713 5154 -410
rect 5418 -1885 5460 -613
rect 5512 -1713 5554 -410
rect 5818 -1885 5860 -613
rect 5912 -1713 5954 -410
rect 6218 -1885 6260 -613
rect 6312 -1713 6354 -410
rect 6618 -1885 6660 -613
rect 6712 -1713 6754 -410
rect 7018 -1885 7060 -613
rect 7112 -1713 7154 -410
rect 7418 -1885 7460 -613
rect 7512 -1713 7554 -410
rect 7818 -1885 7860 -613
rect 7912 -1713 7954 -410
rect 8218 -1885 8260 -613
rect 8312 -1713 8354 -410
rect 8618 -1885 8660 -613
rect 8712 -1713 8754 -410
rect 9018 -1885 9060 -613
rect 9112 -1713 9154 -410
rect 9418 -1885 9460 -613
rect 9512 -1713 9554 -410
rect 9818 -1885 9860 -613
rect 3818 -1890 9860 -1885
rect 3818 -1918 10047 -1890
rect 7784 -2065 8276 -2034
rect 7784 -2075 7825 -2065
rect 7449 -2076 7825 -2075
rect 5555 -2077 7825 -2076
rect 3391 -2106 7825 -2077
rect 3391 -2110 6233 -2106
rect 3391 -3413 3433 -2110
rect 3697 -3585 3739 -2313
rect 3791 -3413 3833 -2110
rect 4097 -3585 4139 -2313
rect 4191 -3413 4233 -2110
rect 4497 -3585 4539 -2313
rect 4591 -3413 4633 -2110
rect 4897 -3585 4939 -2313
rect 4991 -3413 5033 -2110
rect 5297 -3585 5339 -2313
rect 5391 -3413 5433 -2110
rect 5697 -3585 5739 -2313
rect 5791 -3413 5833 -2110
rect 6097 -3585 6139 -2313
rect 6191 -3413 6233 -2110
rect 7350 -2146 7825 -2106
rect 6497 -3585 6539 -2313
rect 7350 -2358 7476 -2146
rect 7784 -2162 7825 -2146
rect 8240 -2162 8276 -2065
rect 9210 -2151 10047 -1918
rect 7784 -2182 8276 -2162
rect 7029 -2398 7789 -2358
rect 9534 -2390 9650 -2151
rect 7029 -2766 7077 -2398
rect 7741 -2719 7789 -2398
rect 8294 -2428 9842 -2390
rect 7741 -2766 7901 -2719
rect 7172 -3252 7235 -2826
rect 7284 -2853 7537 -2807
rect 7836 -2835 7901 -2766
rect 8294 -2795 8336 -2428
rect 7836 -2882 8426 -2835
rect 8600 -2990 8650 -2595
rect 8694 -2795 8736 -2428
rect 8995 -2795 9136 -2736
rect 9400 -2795 9442 -2428
rect 9043 -2990 9093 -2795
rect 9486 -2990 9536 -2595
rect 9800 -2795 9842 -2428
rect 8600 -3029 9536 -2990
rect 8865 -3118 8895 -3029
rect 9235 -3118 9258 -3029
rect 8865 -3132 9258 -3118
rect 8224 -3188 8526 -3157
rect 6725 -3306 7565 -3252
rect 6725 -3407 6799 -3306
rect 6725 -3505 6767 -3407
rect 7501 -3501 7565 -3306
rect 7309 -3505 7565 -3501
rect 6725 -3537 7565 -3505
rect 8224 -3503 8261 -3188
rect 8486 -3503 8526 -3188
rect 8224 -3540 8526 -3503
rect 3697 -3616 6539 -3585
rect 3697 -3618 4192 -3616
rect 4134 -3715 4192 -3618
rect 5698 -3618 6539 -3616
rect 5698 -3715 5736 -3618
rect 4134 -3737 5736 -3715
<< via1 >>
rect 6799 -3407 7501 -3306
rect 6799 -3501 7309 -3407
rect 7309 -3501 7501 -3407
<< metal2 >>
rect 6725 -3306 7565 -3252
rect 6725 -3501 6799 -3306
rect 7501 -3501 7565 -3306
rect 6725 -3537 7565 -3501
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_0
timestamp 1697035654
transform 1 0 4886 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_1
timestamp 1697035654
transform 1 0 3686 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_2
timestamp 1697035654
transform 1 0 4086 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_3
timestamp 1697035654
transform 1 0 4486 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_4
timestamp 1697035654
transform 1 0 6086 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_5
timestamp 1697035654
transform 1 0 5286 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_6
timestamp 1697035654
transform 1 0 5686 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_7
timestamp 1697035654
transform 1 0 6886 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_8
timestamp 1697035654
transform 1 0 6486 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_16
timestamp 1697035654
transform 1 0 3565 0 -1 -2863
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_17
timestamp 1697035654
transform 1 0 3965 0 -1 -2863
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_18
timestamp 1697035654
transform 1 0 4365 0 -1 -2863
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_19
timestamp 1697035654
transform 1 0 4765 0 -1 -2863
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_20
timestamp 1697035654
transform 1 0 5165 0 -1 -2863
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_21
timestamp 1697035654
transform 1 0 5565 0 -1 -2863
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_22
timestamp 1697035654
transform 1 0 5965 0 -1 -2863
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_23
timestamp 1697035654
transform 1 0 6365 0 -1 -2863
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_25
timestamp 1697035654
transform 1 0 9686 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_26
timestamp 1697035654
transform 1 0 9286 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_27
timestamp 1697035654
transform 1 0 8886 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_28
timestamp 1697035654
transform 1 0 8486 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_29
timestamp 1697035654
transform 1 0 8086 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_30
timestamp 1697035654
transform 1 0 7686 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__nfet_01v8_lvt_P9XYHJ  sky130_fd_pr__nfet_01v8_lvt_P9XYHJ_31
timestamp 1697035654
transform 1 0 7286 0 -1 -1163
box -138 -638 138 638
use sky130_fd_pr__pfet_01v8_lvt_G2G9KE  sky130_fd_pr__pfet_01v8_lvt_G2G9KE_0
timestamp 1697034391
transform 1 0 7209 0 -1 -2666
box -174 -200 174 200
use sky130_fd_pr__pfet_01v8_lvt_G2G9KE  sky130_fd_pr__pfet_01v8_lvt_G2G9KE_1
timestamp 1697034391
transform 1 0 7609 0 -1 -2666
box -174 -200 174 200
use sky130_fd_pr__pfet_01v8_lvt_G2G9KE  sky130_fd_pr__pfet_01v8_lvt_G2G9KE_2
timestamp 1697034391
transform 1 0 9668 0 -1 -2695
box -174 -200 174 200
use sky130_fd_pr__pfet_01v8_lvt_G2G9KE  sky130_fd_pr__pfet_01v8_lvt_G2G9KE_3
timestamp 1697034391
transform 1 0 8468 0 -1 -2695
box -174 -200 174 200
use sky130_fd_pr__pfet_01v8_lvt_G2G9KE  sky130_fd_pr__pfet_01v8_lvt_G2G9KE_4
timestamp 1697034391
transform 1 0 8868 0 -1 -2695
box -174 -200 174 200
use sky130_fd_pr__pfet_01v8_lvt_G2G9KE  sky130_fd_pr__pfet_01v8_lvt_G2G9KE_5
timestamp 1697034391
transform 1 0 9268 0 -1 -2695
box -174 -200 174 200
<< labels >>
flabel metal1 9709 -2080 9837 -1976 0 FreeSans 1600 0 0 0 OUT
flabel metal2 7410 -3390 7538 -3286 0 FreeSans 1600 0 0 0 IN
flabel viali 8315 -3415 8443 -3311 0 FreeSans 1600 0 0 0 DD
flabel locali 3197 -3727 3325 -3623 0 FreeSans 1600 0 0 0 SS
<< end >>

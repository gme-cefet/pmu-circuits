magic
tech sky130A
magscale 1 2
timestamp 1698860844
<< nwell >>
rect 106133 277914 107804 279258
rect 106272 276894 107744 277360
rect 106670 274677 109883 275970
rect 114419 272669 115786 280999
rect 120201 279136 121769 280849
rect 122142 280643 123674 280644
rect 120201 273034 121764 279136
rect 122133 278930 123674 280643
rect 122218 277151 124406 278518
rect 122242 276273 124028 276887
rect 122247 275515 124993 276007
rect 109052 270485 109897 272638
rect 112237 270724 115567 271722
rect 120201 268958 123590 273034
rect 120201 268942 121884 268958
<< pwell >>
rect 109581 276507 110259 279221
rect 122756 274452 124148 275072
<< nmos >>
rect 106981 271807 107191 271971
<< pmos >>
rect 106951 274935 107129 275713
rect 107451 274935 107629 275713
rect 107951 274935 108129 275713
rect 108451 274935 108629 275713
rect 108951 274935 109129 275713
rect 109451 274935 109629 275713
rect 122414 277792 123290 278266
rect 122466 275711 122866 275811
rect 123102 275711 123502 275811
rect 123738 275711 124138 275811
rect 124374 275711 124774 275811
<< pmoslvt >>
rect 106368 278757 107582 279011
rect 106368 278157 107582 278411
rect 106491 277090 107525 277164
rect 109440 270706 109510 272426
rect 114657 280403 114857 280803
rect 114657 279957 114857 280117
rect 114657 279549 114857 279709
rect 115348 280403 115548 280803
rect 115348 279957 115548 280117
rect 115348 279549 115548 279709
rect 114657 278737 114857 279137
rect 114657 278291 114857 278451
rect 114657 277883 114857 278043
rect 115348 278737 115548 279137
rect 115348 278291 115548 278451
rect 115348 277883 115548 278043
rect 114657 277071 114857 277471
rect 114657 276625 114857 276785
rect 114657 276217 114857 276377
rect 115348 277071 115548 277471
rect 115348 276625 115548 276785
rect 115348 276217 115548 276377
rect 114657 275405 114857 275805
rect 114657 274959 114857 275119
rect 114657 274551 114857 274711
rect 115348 275405 115548 275805
rect 115348 274959 115548 275119
rect 115348 274551 115548 274711
rect 114657 273739 114857 274139
rect 114657 273293 114857 273453
rect 114657 272885 114857 273045
rect 115348 273739 115548 274139
rect 115348 273293 115548 273453
rect 115348 272885 115548 273045
rect 112578 271106 112738 271306
rect 112978 271106 113138 271306
rect 113378 271106 113538 271306
rect 113778 271106 113938 271306
rect 114637 271077 114797 271277
rect 115037 271077 115197 271277
rect 120429 280537 120829 280637
rect 121129 280537 121529 280637
rect 120429 279753 120829 280253
rect 121129 279753 121529 280253
rect 120429 278969 120829 279469
rect 121129 278969 121529 279469
rect 120429 278185 120829 278685
rect 121129 278185 121529 278685
rect 120429 277401 120829 277901
rect 121129 277401 121529 277901
rect 120429 276617 120829 277117
rect 121129 276617 121529 277117
rect 120429 275833 120829 276333
rect 121129 275833 121529 276333
rect 120429 275049 120829 275549
rect 121129 275049 121529 275549
rect 120429 274265 120829 274765
rect 121129 274265 121529 274765
rect 120429 273481 120829 273981
rect 121129 273481 121529 273981
rect 120429 272697 120829 273197
rect 121129 272697 121529 273197
rect 120429 271913 120829 272413
rect 121129 271913 121529 272413
rect 120429 271129 120829 271629
rect 121129 271129 121529 271629
rect 120429 270345 120829 270845
rect 121129 270345 121529 270845
rect 120429 269561 120829 270061
rect 121129 269561 121529 270061
rect 120429 269177 120829 269277
rect 121129 269177 121529 269277
rect 122356 279923 122756 280423
rect 123056 279923 123456 280423
rect 122356 279139 122756 279639
rect 123056 279139 123456 279639
rect 122416 277400 123216 277500
rect 123656 277394 124210 278080
rect 122438 276492 123832 276668
rect 122125 272713 122525 272813
rect 122825 272713 123225 272813
rect 122125 271929 122525 272429
rect 122825 271929 123225 272429
rect 122125 271145 122525 271645
rect 122825 271145 123225 271645
rect 122125 270361 122525 270861
rect 122825 270361 123225 270861
rect 122125 269577 122525 270077
rect 122825 269577 123225 270077
rect 122125 269193 122525 269293
rect 122825 269193 123225 269293
<< nmoslvt >>
rect 106357 279793 106489 280813
rect 106757 279793 106889 280813
rect 107157 279793 107289 280813
rect 107557 279793 107689 280813
rect 107957 279793 108089 280813
rect 108357 279793 108489 280813
rect 108757 279793 108889 280813
rect 109157 279793 109289 280813
rect 109557 279793 109689 280813
rect 109957 279793 110089 280813
rect 109777 277973 110063 279011
rect 109777 276717 110063 277755
rect 107459 271735 108079 272079
rect 107173 271311 108373 271489
rect 107173 270941 108373 271119
rect 111524 280660 112624 280820
rect 112970 280628 114070 280828
rect 111524 280300 112624 280460
rect 112970 280204 114070 280404
rect 111524 279940 112624 280100
rect 113000 279922 114100 280002
rect 111524 279580 112624 279740
rect 113000 279624 114100 279704
rect 116135 280628 117235 280828
rect 117581 280660 118681 280820
rect 116135 280204 117235 280404
rect 117581 280300 118681 280460
rect 116105 279922 117205 280002
rect 117581 279940 118681 280100
rect 116105 279624 117205 279704
rect 117581 279580 118681 279740
rect 111524 278994 112624 279154
rect 112970 278962 114070 279162
rect 111524 278634 112624 278794
rect 112970 278538 114070 278738
rect 111524 278274 112624 278434
rect 113000 278256 114100 278336
rect 111524 277914 112624 278074
rect 113000 277958 114100 278038
rect 116135 278962 117235 279162
rect 117581 278994 118681 279154
rect 116135 278538 117235 278738
rect 117581 278634 118681 278794
rect 116105 278256 117205 278336
rect 117581 278274 118681 278434
rect 116105 277958 117205 278038
rect 117581 277914 118681 278074
rect 111524 277328 112624 277488
rect 112970 277296 114070 277496
rect 111524 276968 112624 277128
rect 112970 276872 114070 277072
rect 111524 276608 112624 276768
rect 113000 276590 114100 276670
rect 111524 276248 112624 276408
rect 113000 276292 114100 276372
rect 116135 277296 117235 277496
rect 117581 277328 118681 277488
rect 116135 276872 117235 277072
rect 117581 276968 118681 277128
rect 116105 276590 117205 276670
rect 117581 276608 118681 276768
rect 116105 276292 117205 276372
rect 117581 276248 118681 276408
rect 111524 275662 112624 275822
rect 112970 275630 114070 275830
rect 111524 275302 112624 275462
rect 112970 275206 114070 275406
rect 111524 274942 112624 275102
rect 113000 274924 114100 275004
rect 111524 274582 112624 274742
rect 113000 274626 114100 274706
rect 116135 275630 117235 275830
rect 117581 275662 118681 275822
rect 116135 275206 117235 275406
rect 117581 275302 118681 275462
rect 116105 274924 117205 275004
rect 117581 274942 118681 275102
rect 116105 274626 117205 274706
rect 117581 274582 118681 274742
rect 111524 273996 112624 274156
rect 112970 273964 114070 274164
rect 111524 273636 112624 273796
rect 112970 273540 114070 273740
rect 111524 273276 112624 273436
rect 113000 273258 114100 273338
rect 111524 272916 112624 273076
rect 113000 272960 114100 273040
rect 116135 273964 117235 274164
rect 117581 273996 118681 274156
rect 116135 273540 117235 273740
rect 117581 273636 118681 273796
rect 116105 273258 117205 273338
rect 117581 273276 118681 273436
rect 116105 272960 117205 273040
rect 117581 272916 118681 273076
rect 115881 270824 116041 271924
rect 116281 270824 116441 271924
rect 116681 270824 116841 271924
rect 117081 270824 117241 271924
rect 117481 270824 117641 271924
rect 117881 270824 118041 271924
rect 118281 270824 118441 271924
rect 118681 270824 118841 271924
rect 112560 269124 112720 270224
rect 112960 269124 113120 270224
rect 113360 269124 113520 270224
rect 113760 269124 113920 270224
rect 114160 269124 114320 270224
rect 114560 269124 114720 270224
rect 114960 269124 115120 270224
rect 115360 269124 115520 270224
rect 115760 269124 115920 270224
rect 116160 269124 116320 270224
rect 116560 269124 116720 270224
rect 116960 269124 117120 270224
rect 117360 269124 117520 270224
rect 117760 269124 117920 270224
rect 118160 269124 118320 270224
rect 118560 269124 118720 270224
rect 122952 274662 123952 274862
rect 122277 273778 122477 274278
rect 122693 273778 122893 274278
rect 123109 273778 123309 274278
rect 123525 273778 123725 274278
rect 123941 273778 124141 274278
rect 124357 273778 124557 274278
rect 124192 272320 124692 272520
rect 124192 271904 124692 272104
rect 124192 271488 124692 271688
rect 124192 271072 124692 271272
rect 124192 270656 124692 270856
rect 124192 270240 124692 270440
rect 124192 269824 124692 270024
rect 124192 269408 124692 269608
<< ndiff >>
rect 106299 280801 106357 280813
rect 106299 279805 106311 280801
rect 106345 279805 106357 280801
rect 106299 279793 106357 279805
rect 106489 280801 106547 280813
rect 106489 279805 106501 280801
rect 106535 279805 106547 280801
rect 106489 279793 106547 279805
rect 106699 280801 106757 280813
rect 106699 279805 106711 280801
rect 106745 279805 106757 280801
rect 106699 279793 106757 279805
rect 106889 280801 106947 280813
rect 106889 279805 106901 280801
rect 106935 279805 106947 280801
rect 106889 279793 106947 279805
rect 107099 280801 107157 280813
rect 107099 279805 107111 280801
rect 107145 279805 107157 280801
rect 107099 279793 107157 279805
rect 107289 280801 107347 280813
rect 107289 279805 107301 280801
rect 107335 279805 107347 280801
rect 107289 279793 107347 279805
rect 107499 280801 107557 280813
rect 107499 279805 107511 280801
rect 107545 279805 107557 280801
rect 107499 279793 107557 279805
rect 107689 280801 107747 280813
rect 107689 279805 107701 280801
rect 107735 279805 107747 280801
rect 107689 279793 107747 279805
rect 107899 280801 107957 280813
rect 107899 279805 107911 280801
rect 107945 279805 107957 280801
rect 107899 279793 107957 279805
rect 108089 280801 108147 280813
rect 108089 279805 108101 280801
rect 108135 279805 108147 280801
rect 108089 279793 108147 279805
rect 108299 280801 108357 280813
rect 108299 279805 108311 280801
rect 108345 279805 108357 280801
rect 108299 279793 108357 279805
rect 108489 280801 108547 280813
rect 108489 279805 108501 280801
rect 108535 279805 108547 280801
rect 108489 279793 108547 279805
rect 108699 280801 108757 280813
rect 108699 279805 108711 280801
rect 108745 279805 108757 280801
rect 108699 279793 108757 279805
rect 108889 280801 108947 280813
rect 108889 279805 108901 280801
rect 108935 279805 108947 280801
rect 108889 279793 108947 279805
rect 109099 280801 109157 280813
rect 109099 279805 109111 280801
rect 109145 279805 109157 280801
rect 109099 279793 109157 279805
rect 109289 280801 109347 280813
rect 109289 279805 109301 280801
rect 109335 279805 109347 280801
rect 109289 279793 109347 279805
rect 109499 280801 109557 280813
rect 109499 279805 109511 280801
rect 109545 279805 109557 280801
rect 109499 279793 109557 279805
rect 109689 280801 109747 280813
rect 109689 279805 109701 280801
rect 109735 279805 109747 280801
rect 109689 279793 109747 279805
rect 109899 280801 109957 280813
rect 109899 279805 109911 280801
rect 109945 279805 109957 280801
rect 109899 279793 109957 279805
rect 110089 280801 110147 280813
rect 110089 279805 110101 280801
rect 110135 279805 110147 280801
rect 110089 279793 110147 279805
rect 109719 278999 109777 279011
rect 109719 277985 109731 278999
rect 109765 277985 109777 278999
rect 109719 277973 109777 277985
rect 110063 278999 110121 279011
rect 110063 277985 110075 278999
rect 110109 277985 110121 278999
rect 110063 277973 110121 277985
rect 109719 277743 109777 277755
rect 109719 276729 109731 277743
rect 109765 276729 109777 277743
rect 109719 276717 109777 276729
rect 110063 277743 110121 277755
rect 110063 276729 110075 277743
rect 110109 276729 110121 277743
rect 110063 276717 110121 276729
rect 107401 272067 107459 272079
rect 106923 271959 106981 271971
rect 106923 271819 106935 271959
rect 106969 271819 106981 271959
rect 106923 271807 106981 271819
rect 107191 271959 107249 271971
rect 107191 271819 107203 271959
rect 107237 271819 107249 271959
rect 107191 271807 107249 271819
rect 107401 271747 107413 272067
rect 107447 271747 107459 272067
rect 107401 271735 107459 271747
rect 108079 272067 108137 272079
rect 108079 271747 108091 272067
rect 108125 271747 108137 272067
rect 108079 271735 108137 271747
rect 107173 271535 108373 271547
rect 107173 271501 107185 271535
rect 108361 271501 108373 271535
rect 107173 271489 108373 271501
rect 107173 271299 108373 271311
rect 107173 271265 107185 271299
rect 108361 271265 108373 271299
rect 107173 271253 108373 271265
rect 107173 271165 108373 271177
rect 107173 271131 107185 271165
rect 108361 271131 108373 271165
rect 107173 271119 108373 271131
rect 107173 270929 108373 270941
rect 107173 270895 107185 270929
rect 108361 270895 108373 270929
rect 107173 270883 108373 270895
rect 111524 280866 112624 280878
rect 111524 280832 111536 280866
rect 112612 280832 112624 280866
rect 111524 280820 112624 280832
rect 112970 280874 114070 280886
rect 112970 280840 112982 280874
rect 114058 280840 114070 280874
rect 112970 280828 114070 280840
rect 111524 280648 112624 280660
rect 111524 280614 111536 280648
rect 112612 280614 112624 280648
rect 111524 280602 112624 280614
rect 112970 280616 114070 280628
rect 112970 280582 112982 280616
rect 114058 280582 114070 280616
rect 112970 280570 114070 280582
rect 111524 280506 112624 280518
rect 111524 280472 111536 280506
rect 112612 280472 112624 280506
rect 111524 280460 112624 280472
rect 112970 280450 114070 280462
rect 112970 280416 112982 280450
rect 114058 280416 114070 280450
rect 112970 280404 114070 280416
rect 111524 280288 112624 280300
rect 111524 280254 111536 280288
rect 112612 280254 112624 280288
rect 111524 280242 112624 280254
rect 112970 280192 114070 280204
rect 112970 280158 112982 280192
rect 114058 280158 114070 280192
rect 111524 280146 112624 280158
rect 112970 280146 114070 280158
rect 111524 280112 111536 280146
rect 112612 280112 112624 280146
rect 111524 280100 112624 280112
rect 113000 280048 114100 280060
rect 113000 280014 113012 280048
rect 114088 280014 114100 280048
rect 113000 280002 114100 280014
rect 111524 279928 112624 279940
rect 111524 279894 111536 279928
rect 112612 279894 112624 279928
rect 111524 279882 112624 279894
rect 113000 279910 114100 279922
rect 113000 279876 113012 279910
rect 114088 279876 114100 279910
rect 113000 279864 114100 279876
rect 111524 279786 112624 279798
rect 111524 279752 111536 279786
rect 112612 279752 112624 279786
rect 111524 279740 112624 279752
rect 113000 279750 114100 279762
rect 113000 279716 113012 279750
rect 114088 279716 114100 279750
rect 113000 279704 114100 279716
rect 113000 279612 114100 279624
rect 111524 279568 112624 279580
rect 111524 279534 111536 279568
rect 112612 279534 112624 279568
rect 113000 279578 113012 279612
rect 114088 279578 114100 279612
rect 113000 279566 114100 279578
rect 111524 279522 112624 279534
rect 116135 280874 117235 280886
rect 116135 280840 116147 280874
rect 117223 280840 117235 280874
rect 116135 280828 117235 280840
rect 117581 280866 118681 280878
rect 117581 280832 117593 280866
rect 118669 280832 118681 280866
rect 117581 280820 118681 280832
rect 117581 280648 118681 280660
rect 116135 280616 117235 280628
rect 116135 280582 116147 280616
rect 117223 280582 117235 280616
rect 117581 280614 117593 280648
rect 118669 280614 118681 280648
rect 117581 280602 118681 280614
rect 116135 280570 117235 280582
rect 117581 280506 118681 280518
rect 117581 280472 117593 280506
rect 118669 280472 118681 280506
rect 116135 280450 117235 280462
rect 117581 280460 118681 280472
rect 116135 280416 116147 280450
rect 117223 280416 117235 280450
rect 116135 280404 117235 280416
rect 117581 280288 118681 280300
rect 117581 280254 117593 280288
rect 118669 280254 118681 280288
rect 117581 280242 118681 280254
rect 116135 280192 117235 280204
rect 116135 280158 116147 280192
rect 117223 280158 117235 280192
rect 116135 280146 117235 280158
rect 117581 280146 118681 280158
rect 117581 280112 117593 280146
rect 118669 280112 118681 280146
rect 117581 280100 118681 280112
rect 116105 280048 117205 280060
rect 116105 280014 116117 280048
rect 117193 280014 117205 280048
rect 116105 280002 117205 280014
rect 117581 279928 118681 279940
rect 116105 279910 117205 279922
rect 116105 279876 116117 279910
rect 117193 279876 117205 279910
rect 117581 279894 117593 279928
rect 118669 279894 118681 279928
rect 117581 279882 118681 279894
rect 116105 279864 117205 279876
rect 117581 279786 118681 279798
rect 116105 279750 117205 279762
rect 116105 279716 116117 279750
rect 117193 279716 117205 279750
rect 117581 279752 117593 279786
rect 118669 279752 118681 279786
rect 117581 279740 118681 279752
rect 116105 279704 117205 279716
rect 116105 279612 117205 279624
rect 116105 279578 116117 279612
rect 117193 279578 117205 279612
rect 116105 279566 117205 279578
rect 117581 279568 118681 279580
rect 117581 279534 117593 279568
rect 118669 279534 118681 279568
rect 117581 279522 118681 279534
rect 111524 279200 112624 279212
rect 111524 279166 111536 279200
rect 112612 279166 112624 279200
rect 111524 279154 112624 279166
rect 112970 279208 114070 279220
rect 112970 279174 112982 279208
rect 114058 279174 114070 279208
rect 112970 279162 114070 279174
rect 111524 278982 112624 278994
rect 111524 278948 111536 278982
rect 112612 278948 112624 278982
rect 111524 278936 112624 278948
rect 112970 278950 114070 278962
rect 112970 278916 112982 278950
rect 114058 278916 114070 278950
rect 112970 278904 114070 278916
rect 111524 278840 112624 278852
rect 111524 278806 111536 278840
rect 112612 278806 112624 278840
rect 111524 278794 112624 278806
rect 112970 278784 114070 278796
rect 112970 278750 112982 278784
rect 114058 278750 114070 278784
rect 112970 278738 114070 278750
rect 111524 278622 112624 278634
rect 111524 278588 111536 278622
rect 112612 278588 112624 278622
rect 111524 278576 112624 278588
rect 112970 278526 114070 278538
rect 112970 278492 112982 278526
rect 114058 278492 114070 278526
rect 111524 278480 112624 278492
rect 112970 278480 114070 278492
rect 111524 278446 111536 278480
rect 112612 278446 112624 278480
rect 111524 278434 112624 278446
rect 113000 278382 114100 278394
rect 113000 278348 113012 278382
rect 114088 278348 114100 278382
rect 113000 278336 114100 278348
rect 111524 278262 112624 278274
rect 111524 278228 111536 278262
rect 112612 278228 112624 278262
rect 111524 278216 112624 278228
rect 113000 278244 114100 278256
rect 113000 278210 113012 278244
rect 114088 278210 114100 278244
rect 113000 278198 114100 278210
rect 111524 278120 112624 278132
rect 111524 278086 111536 278120
rect 112612 278086 112624 278120
rect 111524 278074 112624 278086
rect 113000 278084 114100 278096
rect 113000 278050 113012 278084
rect 114088 278050 114100 278084
rect 113000 278038 114100 278050
rect 113000 277946 114100 277958
rect 111524 277902 112624 277914
rect 111524 277868 111536 277902
rect 112612 277868 112624 277902
rect 113000 277912 113012 277946
rect 114088 277912 114100 277946
rect 113000 277900 114100 277912
rect 111524 277856 112624 277868
rect 116135 279208 117235 279220
rect 116135 279174 116147 279208
rect 117223 279174 117235 279208
rect 116135 279162 117235 279174
rect 117581 279200 118681 279212
rect 117581 279166 117593 279200
rect 118669 279166 118681 279200
rect 117581 279154 118681 279166
rect 117581 278982 118681 278994
rect 116135 278950 117235 278962
rect 116135 278916 116147 278950
rect 117223 278916 117235 278950
rect 117581 278948 117593 278982
rect 118669 278948 118681 278982
rect 117581 278936 118681 278948
rect 116135 278904 117235 278916
rect 117581 278840 118681 278852
rect 117581 278806 117593 278840
rect 118669 278806 118681 278840
rect 116135 278784 117235 278796
rect 117581 278794 118681 278806
rect 116135 278750 116147 278784
rect 117223 278750 117235 278784
rect 116135 278738 117235 278750
rect 117581 278622 118681 278634
rect 117581 278588 117593 278622
rect 118669 278588 118681 278622
rect 117581 278576 118681 278588
rect 116135 278526 117235 278538
rect 116135 278492 116147 278526
rect 117223 278492 117235 278526
rect 116135 278480 117235 278492
rect 117581 278480 118681 278492
rect 117581 278446 117593 278480
rect 118669 278446 118681 278480
rect 117581 278434 118681 278446
rect 116105 278382 117205 278394
rect 116105 278348 116117 278382
rect 117193 278348 117205 278382
rect 116105 278336 117205 278348
rect 117581 278262 118681 278274
rect 116105 278244 117205 278256
rect 116105 278210 116117 278244
rect 117193 278210 117205 278244
rect 117581 278228 117593 278262
rect 118669 278228 118681 278262
rect 117581 278216 118681 278228
rect 116105 278198 117205 278210
rect 117581 278120 118681 278132
rect 116105 278084 117205 278096
rect 116105 278050 116117 278084
rect 117193 278050 117205 278084
rect 117581 278086 117593 278120
rect 118669 278086 118681 278120
rect 117581 278074 118681 278086
rect 116105 278038 117205 278050
rect 116105 277946 117205 277958
rect 116105 277912 116117 277946
rect 117193 277912 117205 277946
rect 116105 277900 117205 277912
rect 117581 277902 118681 277914
rect 117581 277868 117593 277902
rect 118669 277868 118681 277902
rect 117581 277856 118681 277868
rect 111524 277534 112624 277546
rect 111524 277500 111536 277534
rect 112612 277500 112624 277534
rect 111524 277488 112624 277500
rect 112970 277542 114070 277554
rect 112970 277508 112982 277542
rect 114058 277508 114070 277542
rect 112970 277496 114070 277508
rect 111524 277316 112624 277328
rect 111524 277282 111536 277316
rect 112612 277282 112624 277316
rect 111524 277270 112624 277282
rect 112970 277284 114070 277296
rect 112970 277250 112982 277284
rect 114058 277250 114070 277284
rect 112970 277238 114070 277250
rect 111524 277174 112624 277186
rect 111524 277140 111536 277174
rect 112612 277140 112624 277174
rect 111524 277128 112624 277140
rect 112970 277118 114070 277130
rect 112970 277084 112982 277118
rect 114058 277084 114070 277118
rect 112970 277072 114070 277084
rect 111524 276956 112624 276968
rect 111524 276922 111536 276956
rect 112612 276922 112624 276956
rect 111524 276910 112624 276922
rect 112970 276860 114070 276872
rect 112970 276826 112982 276860
rect 114058 276826 114070 276860
rect 111524 276814 112624 276826
rect 112970 276814 114070 276826
rect 111524 276780 111536 276814
rect 112612 276780 112624 276814
rect 111524 276768 112624 276780
rect 113000 276716 114100 276728
rect 113000 276682 113012 276716
rect 114088 276682 114100 276716
rect 113000 276670 114100 276682
rect 111524 276596 112624 276608
rect 111524 276562 111536 276596
rect 112612 276562 112624 276596
rect 111524 276550 112624 276562
rect 113000 276578 114100 276590
rect 113000 276544 113012 276578
rect 114088 276544 114100 276578
rect 113000 276532 114100 276544
rect 111524 276454 112624 276466
rect 111524 276420 111536 276454
rect 112612 276420 112624 276454
rect 111524 276408 112624 276420
rect 113000 276418 114100 276430
rect 113000 276384 113012 276418
rect 114088 276384 114100 276418
rect 113000 276372 114100 276384
rect 113000 276280 114100 276292
rect 111524 276236 112624 276248
rect 111524 276202 111536 276236
rect 112612 276202 112624 276236
rect 113000 276246 113012 276280
rect 114088 276246 114100 276280
rect 113000 276234 114100 276246
rect 111524 276190 112624 276202
rect 116135 277542 117235 277554
rect 116135 277508 116147 277542
rect 117223 277508 117235 277542
rect 116135 277496 117235 277508
rect 117581 277534 118681 277546
rect 117581 277500 117593 277534
rect 118669 277500 118681 277534
rect 117581 277488 118681 277500
rect 117581 277316 118681 277328
rect 116135 277284 117235 277296
rect 116135 277250 116147 277284
rect 117223 277250 117235 277284
rect 117581 277282 117593 277316
rect 118669 277282 118681 277316
rect 117581 277270 118681 277282
rect 116135 277238 117235 277250
rect 117581 277174 118681 277186
rect 117581 277140 117593 277174
rect 118669 277140 118681 277174
rect 116135 277118 117235 277130
rect 117581 277128 118681 277140
rect 116135 277084 116147 277118
rect 117223 277084 117235 277118
rect 116135 277072 117235 277084
rect 117581 276956 118681 276968
rect 117581 276922 117593 276956
rect 118669 276922 118681 276956
rect 117581 276910 118681 276922
rect 116135 276860 117235 276872
rect 116135 276826 116147 276860
rect 117223 276826 117235 276860
rect 116135 276814 117235 276826
rect 117581 276814 118681 276826
rect 117581 276780 117593 276814
rect 118669 276780 118681 276814
rect 117581 276768 118681 276780
rect 116105 276716 117205 276728
rect 116105 276682 116117 276716
rect 117193 276682 117205 276716
rect 116105 276670 117205 276682
rect 117581 276596 118681 276608
rect 116105 276578 117205 276590
rect 116105 276544 116117 276578
rect 117193 276544 117205 276578
rect 117581 276562 117593 276596
rect 118669 276562 118681 276596
rect 117581 276550 118681 276562
rect 116105 276532 117205 276544
rect 117581 276454 118681 276466
rect 116105 276418 117205 276430
rect 116105 276384 116117 276418
rect 117193 276384 117205 276418
rect 117581 276420 117593 276454
rect 118669 276420 118681 276454
rect 117581 276408 118681 276420
rect 116105 276372 117205 276384
rect 116105 276280 117205 276292
rect 116105 276246 116117 276280
rect 117193 276246 117205 276280
rect 116105 276234 117205 276246
rect 117581 276236 118681 276248
rect 117581 276202 117593 276236
rect 118669 276202 118681 276236
rect 117581 276190 118681 276202
rect 111524 275868 112624 275880
rect 111524 275834 111536 275868
rect 112612 275834 112624 275868
rect 111524 275822 112624 275834
rect 112970 275876 114070 275888
rect 112970 275842 112982 275876
rect 114058 275842 114070 275876
rect 112970 275830 114070 275842
rect 111524 275650 112624 275662
rect 111524 275616 111536 275650
rect 112612 275616 112624 275650
rect 111524 275604 112624 275616
rect 112970 275618 114070 275630
rect 112970 275584 112982 275618
rect 114058 275584 114070 275618
rect 112970 275572 114070 275584
rect 111524 275508 112624 275520
rect 111524 275474 111536 275508
rect 112612 275474 112624 275508
rect 111524 275462 112624 275474
rect 112970 275452 114070 275464
rect 112970 275418 112982 275452
rect 114058 275418 114070 275452
rect 112970 275406 114070 275418
rect 111524 275290 112624 275302
rect 111524 275256 111536 275290
rect 112612 275256 112624 275290
rect 111524 275244 112624 275256
rect 112970 275194 114070 275206
rect 112970 275160 112982 275194
rect 114058 275160 114070 275194
rect 111524 275148 112624 275160
rect 112970 275148 114070 275160
rect 111524 275114 111536 275148
rect 112612 275114 112624 275148
rect 111524 275102 112624 275114
rect 113000 275050 114100 275062
rect 113000 275016 113012 275050
rect 114088 275016 114100 275050
rect 113000 275004 114100 275016
rect 111524 274930 112624 274942
rect 111524 274896 111536 274930
rect 112612 274896 112624 274930
rect 111524 274884 112624 274896
rect 113000 274912 114100 274924
rect 113000 274878 113012 274912
rect 114088 274878 114100 274912
rect 113000 274866 114100 274878
rect 111524 274788 112624 274800
rect 111524 274754 111536 274788
rect 112612 274754 112624 274788
rect 111524 274742 112624 274754
rect 113000 274752 114100 274764
rect 113000 274718 113012 274752
rect 114088 274718 114100 274752
rect 113000 274706 114100 274718
rect 113000 274614 114100 274626
rect 111524 274570 112624 274582
rect 111524 274536 111536 274570
rect 112612 274536 112624 274570
rect 113000 274580 113012 274614
rect 114088 274580 114100 274614
rect 113000 274568 114100 274580
rect 111524 274524 112624 274536
rect 116135 275876 117235 275888
rect 116135 275842 116147 275876
rect 117223 275842 117235 275876
rect 116135 275830 117235 275842
rect 117581 275868 118681 275880
rect 117581 275834 117593 275868
rect 118669 275834 118681 275868
rect 117581 275822 118681 275834
rect 117581 275650 118681 275662
rect 116135 275618 117235 275630
rect 116135 275584 116147 275618
rect 117223 275584 117235 275618
rect 117581 275616 117593 275650
rect 118669 275616 118681 275650
rect 117581 275604 118681 275616
rect 116135 275572 117235 275584
rect 117581 275508 118681 275520
rect 117581 275474 117593 275508
rect 118669 275474 118681 275508
rect 116135 275452 117235 275464
rect 117581 275462 118681 275474
rect 116135 275418 116147 275452
rect 117223 275418 117235 275452
rect 116135 275406 117235 275418
rect 117581 275290 118681 275302
rect 117581 275256 117593 275290
rect 118669 275256 118681 275290
rect 117581 275244 118681 275256
rect 116135 275194 117235 275206
rect 116135 275160 116147 275194
rect 117223 275160 117235 275194
rect 116135 275148 117235 275160
rect 117581 275148 118681 275160
rect 117581 275114 117593 275148
rect 118669 275114 118681 275148
rect 117581 275102 118681 275114
rect 116105 275050 117205 275062
rect 116105 275016 116117 275050
rect 117193 275016 117205 275050
rect 116105 275004 117205 275016
rect 117581 274930 118681 274942
rect 116105 274912 117205 274924
rect 116105 274878 116117 274912
rect 117193 274878 117205 274912
rect 117581 274896 117593 274930
rect 118669 274896 118681 274930
rect 117581 274884 118681 274896
rect 116105 274866 117205 274878
rect 117581 274788 118681 274800
rect 116105 274752 117205 274764
rect 116105 274718 116117 274752
rect 117193 274718 117205 274752
rect 117581 274754 117593 274788
rect 118669 274754 118681 274788
rect 117581 274742 118681 274754
rect 116105 274706 117205 274718
rect 116105 274614 117205 274626
rect 116105 274580 116117 274614
rect 117193 274580 117205 274614
rect 116105 274568 117205 274580
rect 117581 274570 118681 274582
rect 117581 274536 117593 274570
rect 118669 274536 118681 274570
rect 117581 274524 118681 274536
rect 111524 274202 112624 274214
rect 111524 274168 111536 274202
rect 112612 274168 112624 274202
rect 111524 274156 112624 274168
rect 112970 274210 114070 274222
rect 112970 274176 112982 274210
rect 114058 274176 114070 274210
rect 112970 274164 114070 274176
rect 111524 273984 112624 273996
rect 111524 273950 111536 273984
rect 112612 273950 112624 273984
rect 111524 273938 112624 273950
rect 112970 273952 114070 273964
rect 112970 273918 112982 273952
rect 114058 273918 114070 273952
rect 112970 273906 114070 273918
rect 111524 273842 112624 273854
rect 111524 273808 111536 273842
rect 112612 273808 112624 273842
rect 111524 273796 112624 273808
rect 112970 273786 114070 273798
rect 112970 273752 112982 273786
rect 114058 273752 114070 273786
rect 112970 273740 114070 273752
rect 111524 273624 112624 273636
rect 111524 273590 111536 273624
rect 112612 273590 112624 273624
rect 111524 273578 112624 273590
rect 112970 273528 114070 273540
rect 112970 273494 112982 273528
rect 114058 273494 114070 273528
rect 111524 273482 112624 273494
rect 112970 273482 114070 273494
rect 111524 273448 111536 273482
rect 112612 273448 112624 273482
rect 111524 273436 112624 273448
rect 113000 273384 114100 273396
rect 113000 273350 113012 273384
rect 114088 273350 114100 273384
rect 113000 273338 114100 273350
rect 111524 273264 112624 273276
rect 111524 273230 111536 273264
rect 112612 273230 112624 273264
rect 111524 273218 112624 273230
rect 113000 273246 114100 273258
rect 113000 273212 113012 273246
rect 114088 273212 114100 273246
rect 113000 273200 114100 273212
rect 111524 273122 112624 273134
rect 111524 273088 111536 273122
rect 112612 273088 112624 273122
rect 111524 273076 112624 273088
rect 113000 273086 114100 273098
rect 113000 273052 113012 273086
rect 114088 273052 114100 273086
rect 113000 273040 114100 273052
rect 113000 272948 114100 272960
rect 111524 272904 112624 272916
rect 111524 272870 111536 272904
rect 112612 272870 112624 272904
rect 113000 272914 113012 272948
rect 114088 272914 114100 272948
rect 113000 272902 114100 272914
rect 111524 272858 112624 272870
rect 116135 274210 117235 274222
rect 116135 274176 116147 274210
rect 117223 274176 117235 274210
rect 116135 274164 117235 274176
rect 117581 274202 118681 274214
rect 117581 274168 117593 274202
rect 118669 274168 118681 274202
rect 117581 274156 118681 274168
rect 117581 273984 118681 273996
rect 116135 273952 117235 273964
rect 116135 273918 116147 273952
rect 117223 273918 117235 273952
rect 117581 273950 117593 273984
rect 118669 273950 118681 273984
rect 117581 273938 118681 273950
rect 116135 273906 117235 273918
rect 117581 273842 118681 273854
rect 117581 273808 117593 273842
rect 118669 273808 118681 273842
rect 116135 273786 117235 273798
rect 117581 273796 118681 273808
rect 116135 273752 116147 273786
rect 117223 273752 117235 273786
rect 116135 273740 117235 273752
rect 117581 273624 118681 273636
rect 117581 273590 117593 273624
rect 118669 273590 118681 273624
rect 117581 273578 118681 273590
rect 116135 273528 117235 273540
rect 116135 273494 116147 273528
rect 117223 273494 117235 273528
rect 116135 273482 117235 273494
rect 117581 273482 118681 273494
rect 117581 273448 117593 273482
rect 118669 273448 118681 273482
rect 117581 273436 118681 273448
rect 116105 273384 117205 273396
rect 116105 273350 116117 273384
rect 117193 273350 117205 273384
rect 116105 273338 117205 273350
rect 117581 273264 118681 273276
rect 116105 273246 117205 273258
rect 116105 273212 116117 273246
rect 117193 273212 117205 273246
rect 117581 273230 117593 273264
rect 118669 273230 118681 273264
rect 117581 273218 118681 273230
rect 116105 273200 117205 273212
rect 117581 273122 118681 273134
rect 116105 273086 117205 273098
rect 116105 273052 116117 273086
rect 117193 273052 117205 273086
rect 117581 273088 117593 273122
rect 118669 273088 118681 273122
rect 117581 273076 118681 273088
rect 116105 273040 117205 273052
rect 116105 272948 117205 272960
rect 116105 272914 116117 272948
rect 117193 272914 117205 272948
rect 116105 272902 117205 272914
rect 117581 272904 118681 272916
rect 117581 272870 117593 272904
rect 118669 272870 118681 272904
rect 117581 272858 118681 272870
rect 115823 271912 115881 271924
rect 115823 270836 115835 271912
rect 115869 270836 115881 271912
rect 115823 270824 115881 270836
rect 116041 271912 116099 271924
rect 116041 270836 116053 271912
rect 116087 270836 116099 271912
rect 116041 270824 116099 270836
rect 116223 271912 116281 271924
rect 116223 270836 116235 271912
rect 116269 270836 116281 271912
rect 116223 270824 116281 270836
rect 116441 271912 116499 271924
rect 116441 270836 116453 271912
rect 116487 270836 116499 271912
rect 116441 270824 116499 270836
rect 116623 271912 116681 271924
rect 116623 270836 116635 271912
rect 116669 270836 116681 271912
rect 116623 270824 116681 270836
rect 116841 271912 116899 271924
rect 116841 270836 116853 271912
rect 116887 270836 116899 271912
rect 116841 270824 116899 270836
rect 117023 271912 117081 271924
rect 117023 270836 117035 271912
rect 117069 270836 117081 271912
rect 117023 270824 117081 270836
rect 117241 271912 117299 271924
rect 117241 270836 117253 271912
rect 117287 270836 117299 271912
rect 117241 270824 117299 270836
rect 117423 271912 117481 271924
rect 117423 270836 117435 271912
rect 117469 270836 117481 271912
rect 117423 270824 117481 270836
rect 117641 271912 117699 271924
rect 117641 270836 117653 271912
rect 117687 270836 117699 271912
rect 117641 270824 117699 270836
rect 117823 271912 117881 271924
rect 117823 270836 117835 271912
rect 117869 270836 117881 271912
rect 117823 270824 117881 270836
rect 118041 271912 118099 271924
rect 118041 270836 118053 271912
rect 118087 270836 118099 271912
rect 118041 270824 118099 270836
rect 118223 271912 118281 271924
rect 118223 270836 118235 271912
rect 118269 270836 118281 271912
rect 118223 270824 118281 270836
rect 118441 271912 118499 271924
rect 118441 270836 118453 271912
rect 118487 270836 118499 271912
rect 118441 270824 118499 270836
rect 118623 271912 118681 271924
rect 118623 270836 118635 271912
rect 118669 270836 118681 271912
rect 118623 270824 118681 270836
rect 118841 271912 118899 271924
rect 118841 270836 118853 271912
rect 118887 270836 118899 271912
rect 118841 270824 118899 270836
rect 112502 270212 112560 270224
rect 112502 269136 112514 270212
rect 112548 269136 112560 270212
rect 112502 269124 112560 269136
rect 112720 270212 112778 270224
rect 112720 269136 112732 270212
rect 112766 269136 112778 270212
rect 112720 269124 112778 269136
rect 112902 270212 112960 270224
rect 112902 269136 112914 270212
rect 112948 269136 112960 270212
rect 112902 269124 112960 269136
rect 113120 270212 113178 270224
rect 113120 269136 113132 270212
rect 113166 269136 113178 270212
rect 113120 269124 113178 269136
rect 113302 270212 113360 270224
rect 113302 269136 113314 270212
rect 113348 269136 113360 270212
rect 113302 269124 113360 269136
rect 113520 270212 113578 270224
rect 113520 269136 113532 270212
rect 113566 269136 113578 270212
rect 113520 269124 113578 269136
rect 113702 270212 113760 270224
rect 113702 269136 113714 270212
rect 113748 269136 113760 270212
rect 113702 269124 113760 269136
rect 113920 270212 113978 270224
rect 113920 269136 113932 270212
rect 113966 269136 113978 270212
rect 113920 269124 113978 269136
rect 114102 270212 114160 270224
rect 114102 269136 114114 270212
rect 114148 269136 114160 270212
rect 114102 269124 114160 269136
rect 114320 270212 114378 270224
rect 114320 269136 114332 270212
rect 114366 269136 114378 270212
rect 114320 269124 114378 269136
rect 114502 270212 114560 270224
rect 114502 269136 114514 270212
rect 114548 269136 114560 270212
rect 114502 269124 114560 269136
rect 114720 270212 114778 270224
rect 114720 269136 114732 270212
rect 114766 269136 114778 270212
rect 114720 269124 114778 269136
rect 114902 270212 114960 270224
rect 114902 269136 114914 270212
rect 114948 269136 114960 270212
rect 114902 269124 114960 269136
rect 115120 270212 115178 270224
rect 115120 269136 115132 270212
rect 115166 269136 115178 270212
rect 115120 269124 115178 269136
rect 115302 270212 115360 270224
rect 115302 269136 115314 270212
rect 115348 269136 115360 270212
rect 115302 269124 115360 269136
rect 115520 270212 115578 270224
rect 115520 269136 115532 270212
rect 115566 269136 115578 270212
rect 115520 269124 115578 269136
rect 115702 270212 115760 270224
rect 115702 269136 115714 270212
rect 115748 269136 115760 270212
rect 115702 269124 115760 269136
rect 115920 270212 115978 270224
rect 115920 269136 115932 270212
rect 115966 269136 115978 270212
rect 115920 269124 115978 269136
rect 116102 270212 116160 270224
rect 116102 269136 116114 270212
rect 116148 269136 116160 270212
rect 116102 269124 116160 269136
rect 116320 270212 116378 270224
rect 116320 269136 116332 270212
rect 116366 269136 116378 270212
rect 116320 269124 116378 269136
rect 116502 270212 116560 270224
rect 116502 269136 116514 270212
rect 116548 269136 116560 270212
rect 116502 269124 116560 269136
rect 116720 270212 116778 270224
rect 116720 269136 116732 270212
rect 116766 269136 116778 270212
rect 116720 269124 116778 269136
rect 116902 270212 116960 270224
rect 116902 269136 116914 270212
rect 116948 269136 116960 270212
rect 116902 269124 116960 269136
rect 117120 270212 117178 270224
rect 117120 269136 117132 270212
rect 117166 269136 117178 270212
rect 117120 269124 117178 269136
rect 117302 270212 117360 270224
rect 117302 269136 117314 270212
rect 117348 269136 117360 270212
rect 117302 269124 117360 269136
rect 117520 270212 117578 270224
rect 117520 269136 117532 270212
rect 117566 269136 117578 270212
rect 117520 269124 117578 269136
rect 117702 270212 117760 270224
rect 117702 269136 117714 270212
rect 117748 269136 117760 270212
rect 117702 269124 117760 269136
rect 117920 270212 117978 270224
rect 117920 269136 117932 270212
rect 117966 269136 117978 270212
rect 117920 269124 117978 269136
rect 118102 270212 118160 270224
rect 118102 269136 118114 270212
rect 118148 269136 118160 270212
rect 118102 269124 118160 269136
rect 118320 270212 118378 270224
rect 118320 269136 118332 270212
rect 118366 269136 118378 270212
rect 118320 269124 118378 269136
rect 118502 270212 118560 270224
rect 118502 269136 118514 270212
rect 118548 269136 118560 270212
rect 118502 269124 118560 269136
rect 118720 270212 118778 270224
rect 118720 269136 118732 270212
rect 118766 269136 118778 270212
rect 118720 269124 118778 269136
rect 122894 274850 122952 274862
rect 122894 274674 122906 274850
rect 122940 274674 122952 274850
rect 122894 274662 122952 274674
rect 123952 274850 124010 274862
rect 123952 274674 123964 274850
rect 123998 274674 124010 274850
rect 123952 274662 124010 274674
rect 122219 274266 122277 274278
rect 122219 273790 122231 274266
rect 122265 273790 122277 274266
rect 122219 273778 122277 273790
rect 122477 274266 122535 274278
rect 122477 273790 122489 274266
rect 122523 273790 122535 274266
rect 122477 273778 122535 273790
rect 122635 274266 122693 274278
rect 122635 273790 122647 274266
rect 122681 273790 122693 274266
rect 122635 273778 122693 273790
rect 122893 274266 122951 274278
rect 122893 273790 122905 274266
rect 122939 273790 122951 274266
rect 122893 273778 122951 273790
rect 123051 274266 123109 274278
rect 123051 273790 123063 274266
rect 123097 273790 123109 274266
rect 123051 273778 123109 273790
rect 123309 274266 123367 274278
rect 123309 273790 123321 274266
rect 123355 273790 123367 274266
rect 123309 273778 123367 273790
rect 123467 274266 123525 274278
rect 123467 273790 123479 274266
rect 123513 273790 123525 274266
rect 123467 273778 123525 273790
rect 123725 274266 123783 274278
rect 123725 273790 123737 274266
rect 123771 273790 123783 274266
rect 123725 273778 123783 273790
rect 123883 274266 123941 274278
rect 123883 273790 123895 274266
rect 123929 273790 123941 274266
rect 123883 273778 123941 273790
rect 124141 274266 124199 274278
rect 124141 273790 124153 274266
rect 124187 273790 124199 274266
rect 124141 273778 124199 273790
rect 124299 274266 124357 274278
rect 124299 273790 124311 274266
rect 124345 273790 124357 274266
rect 124299 273778 124357 273790
rect 124557 274266 124615 274278
rect 124557 273790 124569 274266
rect 124603 273790 124615 274266
rect 124557 273778 124615 273790
rect 124192 272566 124692 272578
rect 124192 272532 124204 272566
rect 124680 272532 124692 272566
rect 124192 272520 124692 272532
rect 124192 272308 124692 272320
rect 124192 272274 124204 272308
rect 124680 272274 124692 272308
rect 124192 272262 124692 272274
rect 124192 272150 124692 272162
rect 124192 272116 124204 272150
rect 124680 272116 124692 272150
rect 124192 272104 124692 272116
rect 124192 271892 124692 271904
rect 124192 271858 124204 271892
rect 124680 271858 124692 271892
rect 124192 271846 124692 271858
rect 124192 271734 124692 271746
rect 124192 271700 124204 271734
rect 124680 271700 124692 271734
rect 124192 271688 124692 271700
rect 124192 271476 124692 271488
rect 124192 271442 124204 271476
rect 124680 271442 124692 271476
rect 124192 271430 124692 271442
rect 124192 271318 124692 271330
rect 124192 271284 124204 271318
rect 124680 271284 124692 271318
rect 124192 271272 124692 271284
rect 124192 271060 124692 271072
rect 124192 271026 124204 271060
rect 124680 271026 124692 271060
rect 124192 271014 124692 271026
rect 124192 270902 124692 270914
rect 124192 270868 124204 270902
rect 124680 270868 124692 270902
rect 124192 270856 124692 270868
rect 124192 270644 124692 270656
rect 124192 270610 124204 270644
rect 124680 270610 124692 270644
rect 124192 270598 124692 270610
rect 124192 270486 124692 270498
rect 124192 270452 124204 270486
rect 124680 270452 124692 270486
rect 124192 270440 124692 270452
rect 124192 270228 124692 270240
rect 124192 270194 124204 270228
rect 124680 270194 124692 270228
rect 124192 270182 124692 270194
rect 124192 270070 124692 270082
rect 124192 270036 124204 270070
rect 124680 270036 124692 270070
rect 124192 270024 124692 270036
rect 124192 269812 124692 269824
rect 124192 269778 124204 269812
rect 124680 269778 124692 269812
rect 124192 269766 124692 269778
rect 124192 269654 124692 269666
rect 124192 269620 124204 269654
rect 124680 269620 124692 269654
rect 124192 269608 124692 269620
rect 124192 269396 124692 269408
rect 124192 269362 124204 269396
rect 124680 269362 124692 269396
rect 124192 269350 124692 269362
<< pdiff >>
rect 106368 279057 107582 279069
rect 106368 279023 106380 279057
rect 107570 279023 107582 279057
rect 106368 279011 107582 279023
rect 106368 278745 107582 278757
rect 106368 278711 106380 278745
rect 107570 278711 107582 278745
rect 106368 278699 107582 278711
rect 106368 278457 107582 278469
rect 106368 278423 106380 278457
rect 107570 278423 107582 278457
rect 106368 278411 107582 278423
rect 106368 278145 107582 278157
rect 106368 278111 106380 278145
rect 107570 278111 107582 278145
rect 106368 278099 107582 278111
rect 106491 277210 107525 277222
rect 106491 277176 106503 277210
rect 107513 277176 107525 277210
rect 106491 277164 107525 277176
rect 106491 277078 107525 277090
rect 106491 277044 106503 277078
rect 107513 277044 107525 277078
rect 106491 277032 107525 277044
rect 106951 275759 107129 275771
rect 106951 275725 106963 275759
rect 107117 275725 107129 275759
rect 106951 275713 107129 275725
rect 107451 275759 107629 275771
rect 107451 275725 107463 275759
rect 107617 275725 107629 275759
rect 107451 275713 107629 275725
rect 107951 275759 108129 275771
rect 107951 275725 107963 275759
rect 108117 275725 108129 275759
rect 107951 275713 108129 275725
rect 108451 275759 108629 275771
rect 108451 275725 108463 275759
rect 108617 275725 108629 275759
rect 108451 275713 108629 275725
rect 108951 275759 109129 275771
rect 108951 275725 108963 275759
rect 109117 275725 109129 275759
rect 108951 275713 109129 275725
rect 109451 275759 109629 275771
rect 109451 275725 109463 275759
rect 109617 275725 109629 275759
rect 109451 275713 109629 275725
rect 106951 274923 107129 274935
rect 106951 274889 106963 274923
rect 107117 274889 107129 274923
rect 106951 274877 107129 274889
rect 107451 274923 107629 274935
rect 107451 274889 107463 274923
rect 107617 274889 107629 274923
rect 107451 274877 107629 274889
rect 107951 274923 108129 274935
rect 107951 274889 107963 274923
rect 108117 274889 108129 274923
rect 107951 274877 108129 274889
rect 108451 274923 108629 274935
rect 108451 274889 108463 274923
rect 108617 274889 108629 274923
rect 108451 274877 108629 274889
rect 108951 274923 109129 274935
rect 108951 274889 108963 274923
rect 109117 274889 109129 274923
rect 108951 274877 109129 274889
rect 109451 274923 109629 274935
rect 109451 274889 109463 274923
rect 109617 274889 109629 274923
rect 109451 274877 109629 274889
rect 109240 272414 109440 272426
rect 109240 270718 109394 272414
rect 109428 270718 109440 272414
rect 109240 270706 109440 270718
rect 109510 272414 109710 272426
rect 109510 270718 109522 272414
rect 109556 270718 109710 272414
rect 109510 270706 109710 270718
rect 114657 280849 114857 280861
rect 114657 280815 114669 280849
rect 114845 280815 114857 280849
rect 114657 280803 114857 280815
rect 114657 280391 114857 280403
rect 114657 280357 114669 280391
rect 114845 280357 114857 280391
rect 114657 280345 114857 280357
rect 114657 280163 114857 280175
rect 114657 280129 114669 280163
rect 114845 280129 114857 280163
rect 114657 280117 114857 280129
rect 114657 279945 114857 279957
rect 114657 279911 114669 279945
rect 114845 279911 114857 279945
rect 114657 279899 114857 279911
rect 114657 279755 114857 279767
rect 114657 279721 114669 279755
rect 114845 279721 114857 279755
rect 114657 279709 114857 279721
rect 114657 279537 114857 279549
rect 114657 279503 114669 279537
rect 114845 279503 114857 279537
rect 114657 279491 114857 279503
rect 115348 280849 115548 280861
rect 115348 280815 115360 280849
rect 115536 280815 115548 280849
rect 115348 280803 115548 280815
rect 115348 280391 115548 280403
rect 115348 280357 115360 280391
rect 115536 280357 115548 280391
rect 115348 280345 115548 280357
rect 115348 280163 115548 280175
rect 115348 280129 115360 280163
rect 115536 280129 115548 280163
rect 115348 280117 115548 280129
rect 115348 279945 115548 279957
rect 115348 279911 115360 279945
rect 115536 279911 115548 279945
rect 115348 279899 115548 279911
rect 115348 279755 115548 279767
rect 115348 279721 115360 279755
rect 115536 279721 115548 279755
rect 115348 279709 115548 279721
rect 115348 279537 115548 279549
rect 115348 279503 115360 279537
rect 115536 279503 115548 279537
rect 115348 279491 115548 279503
rect 114657 279183 114857 279195
rect 114657 279149 114669 279183
rect 114845 279149 114857 279183
rect 114657 279137 114857 279149
rect 114657 278725 114857 278737
rect 114657 278691 114669 278725
rect 114845 278691 114857 278725
rect 114657 278679 114857 278691
rect 114657 278497 114857 278509
rect 114657 278463 114669 278497
rect 114845 278463 114857 278497
rect 114657 278451 114857 278463
rect 114657 278279 114857 278291
rect 114657 278245 114669 278279
rect 114845 278245 114857 278279
rect 114657 278233 114857 278245
rect 114657 278089 114857 278101
rect 114657 278055 114669 278089
rect 114845 278055 114857 278089
rect 114657 278043 114857 278055
rect 114657 277871 114857 277883
rect 114657 277837 114669 277871
rect 114845 277837 114857 277871
rect 114657 277825 114857 277837
rect 115348 279183 115548 279195
rect 115348 279149 115360 279183
rect 115536 279149 115548 279183
rect 115348 279137 115548 279149
rect 115348 278725 115548 278737
rect 115348 278691 115360 278725
rect 115536 278691 115548 278725
rect 115348 278679 115548 278691
rect 115348 278497 115548 278509
rect 115348 278463 115360 278497
rect 115536 278463 115548 278497
rect 115348 278451 115548 278463
rect 115348 278279 115548 278291
rect 115348 278245 115360 278279
rect 115536 278245 115548 278279
rect 115348 278233 115548 278245
rect 115348 278089 115548 278101
rect 115348 278055 115360 278089
rect 115536 278055 115548 278089
rect 115348 278043 115548 278055
rect 115348 277871 115548 277883
rect 115348 277837 115360 277871
rect 115536 277837 115548 277871
rect 115348 277825 115548 277837
rect 114657 277517 114857 277529
rect 114657 277483 114669 277517
rect 114845 277483 114857 277517
rect 114657 277471 114857 277483
rect 114657 277059 114857 277071
rect 114657 277025 114669 277059
rect 114845 277025 114857 277059
rect 114657 277013 114857 277025
rect 114657 276831 114857 276843
rect 114657 276797 114669 276831
rect 114845 276797 114857 276831
rect 114657 276785 114857 276797
rect 114657 276613 114857 276625
rect 114657 276579 114669 276613
rect 114845 276579 114857 276613
rect 114657 276567 114857 276579
rect 114657 276423 114857 276435
rect 114657 276389 114669 276423
rect 114845 276389 114857 276423
rect 114657 276377 114857 276389
rect 114657 276205 114857 276217
rect 114657 276171 114669 276205
rect 114845 276171 114857 276205
rect 114657 276159 114857 276171
rect 115348 277517 115548 277529
rect 115348 277483 115360 277517
rect 115536 277483 115548 277517
rect 115348 277471 115548 277483
rect 115348 277059 115548 277071
rect 115348 277025 115360 277059
rect 115536 277025 115548 277059
rect 115348 277013 115548 277025
rect 115348 276831 115548 276843
rect 115348 276797 115360 276831
rect 115536 276797 115548 276831
rect 115348 276785 115548 276797
rect 115348 276613 115548 276625
rect 115348 276579 115360 276613
rect 115536 276579 115548 276613
rect 115348 276567 115548 276579
rect 115348 276423 115548 276435
rect 115348 276389 115360 276423
rect 115536 276389 115548 276423
rect 115348 276377 115548 276389
rect 115348 276205 115548 276217
rect 115348 276171 115360 276205
rect 115536 276171 115548 276205
rect 115348 276159 115548 276171
rect 114657 275851 114857 275863
rect 114657 275817 114669 275851
rect 114845 275817 114857 275851
rect 114657 275805 114857 275817
rect 114657 275393 114857 275405
rect 114657 275359 114669 275393
rect 114845 275359 114857 275393
rect 114657 275347 114857 275359
rect 114657 275165 114857 275177
rect 114657 275131 114669 275165
rect 114845 275131 114857 275165
rect 114657 275119 114857 275131
rect 114657 274947 114857 274959
rect 114657 274913 114669 274947
rect 114845 274913 114857 274947
rect 114657 274901 114857 274913
rect 114657 274757 114857 274769
rect 114657 274723 114669 274757
rect 114845 274723 114857 274757
rect 114657 274711 114857 274723
rect 114657 274539 114857 274551
rect 114657 274505 114669 274539
rect 114845 274505 114857 274539
rect 114657 274493 114857 274505
rect 115348 275851 115548 275863
rect 115348 275817 115360 275851
rect 115536 275817 115548 275851
rect 115348 275805 115548 275817
rect 115348 275393 115548 275405
rect 115348 275359 115360 275393
rect 115536 275359 115548 275393
rect 115348 275347 115548 275359
rect 115348 275165 115548 275177
rect 115348 275131 115360 275165
rect 115536 275131 115548 275165
rect 115348 275119 115548 275131
rect 115348 274947 115548 274959
rect 115348 274913 115360 274947
rect 115536 274913 115548 274947
rect 115348 274901 115548 274913
rect 115348 274757 115548 274769
rect 115348 274723 115360 274757
rect 115536 274723 115548 274757
rect 115348 274711 115548 274723
rect 115348 274539 115548 274551
rect 115348 274505 115360 274539
rect 115536 274505 115548 274539
rect 115348 274493 115548 274505
rect 114657 274185 114857 274197
rect 114657 274151 114669 274185
rect 114845 274151 114857 274185
rect 114657 274139 114857 274151
rect 114657 273727 114857 273739
rect 114657 273693 114669 273727
rect 114845 273693 114857 273727
rect 114657 273681 114857 273693
rect 114657 273499 114857 273511
rect 114657 273465 114669 273499
rect 114845 273465 114857 273499
rect 114657 273453 114857 273465
rect 114657 273281 114857 273293
rect 114657 273247 114669 273281
rect 114845 273247 114857 273281
rect 114657 273235 114857 273247
rect 114657 273091 114857 273103
rect 114657 273057 114669 273091
rect 114845 273057 114857 273091
rect 114657 273045 114857 273057
rect 114657 272873 114857 272885
rect 114657 272839 114669 272873
rect 114845 272839 114857 272873
rect 114657 272827 114857 272839
rect 115348 274185 115548 274197
rect 115348 274151 115360 274185
rect 115536 274151 115548 274185
rect 115348 274139 115548 274151
rect 115348 273727 115548 273739
rect 115348 273693 115360 273727
rect 115536 273693 115548 273727
rect 115348 273681 115548 273693
rect 115348 273499 115548 273511
rect 115348 273465 115360 273499
rect 115536 273465 115548 273499
rect 115348 273453 115548 273465
rect 115348 273281 115548 273293
rect 115348 273247 115360 273281
rect 115536 273247 115548 273281
rect 115348 273235 115548 273247
rect 115348 273091 115548 273103
rect 115348 273057 115360 273091
rect 115536 273057 115548 273091
rect 115348 273045 115548 273057
rect 115348 272873 115548 272885
rect 115348 272839 115360 272873
rect 115536 272839 115548 272873
rect 115348 272827 115548 272839
rect 112520 271294 112578 271306
rect 112520 271118 112532 271294
rect 112566 271118 112578 271294
rect 112520 271106 112578 271118
rect 112738 271294 112796 271306
rect 112738 271118 112750 271294
rect 112784 271118 112796 271294
rect 112738 271106 112796 271118
rect 112920 271294 112978 271306
rect 112920 271118 112932 271294
rect 112966 271118 112978 271294
rect 112920 271106 112978 271118
rect 113138 271294 113196 271306
rect 113138 271118 113150 271294
rect 113184 271118 113196 271294
rect 113138 271106 113196 271118
rect 113320 271294 113378 271306
rect 113320 271118 113332 271294
rect 113366 271118 113378 271294
rect 113320 271106 113378 271118
rect 113538 271294 113596 271306
rect 113538 271118 113550 271294
rect 113584 271118 113596 271294
rect 113538 271106 113596 271118
rect 113720 271294 113778 271306
rect 113720 271118 113732 271294
rect 113766 271118 113778 271294
rect 113720 271106 113778 271118
rect 113938 271294 113996 271306
rect 113938 271118 113950 271294
rect 113984 271118 113996 271294
rect 113938 271106 113996 271118
rect 114579 271265 114637 271277
rect 114579 271089 114591 271265
rect 114625 271089 114637 271265
rect 114579 271077 114637 271089
rect 114797 271265 114855 271277
rect 114797 271089 114809 271265
rect 114843 271089 114855 271265
rect 114797 271077 114855 271089
rect 114979 271265 115037 271277
rect 114979 271089 114991 271265
rect 115025 271089 115037 271265
rect 114979 271077 115037 271089
rect 115197 271265 115255 271277
rect 115197 271089 115209 271265
rect 115243 271089 115255 271265
rect 115197 271077 115255 271089
rect 120371 280625 120429 280637
rect 120371 280549 120383 280625
rect 120417 280549 120429 280625
rect 120371 280537 120429 280549
rect 120829 280625 120887 280637
rect 120829 280549 120841 280625
rect 120875 280549 120887 280625
rect 120829 280537 120887 280549
rect 121071 280625 121129 280637
rect 121071 280549 121083 280625
rect 121117 280549 121129 280625
rect 121071 280537 121129 280549
rect 121529 280625 121587 280637
rect 121529 280549 121541 280625
rect 121575 280549 121587 280625
rect 121529 280537 121587 280549
rect 120371 280241 120429 280253
rect 120371 279765 120383 280241
rect 120417 279765 120429 280241
rect 120371 279753 120429 279765
rect 120829 280241 120887 280253
rect 120829 279765 120841 280241
rect 120875 279765 120887 280241
rect 120829 279753 120887 279765
rect 121071 280241 121129 280253
rect 121071 279765 121083 280241
rect 121117 279765 121129 280241
rect 121071 279753 121129 279765
rect 121529 280241 121587 280253
rect 121529 279765 121541 280241
rect 121575 279765 121587 280241
rect 121529 279753 121587 279765
rect 120371 279457 120429 279469
rect 120371 278981 120383 279457
rect 120417 278981 120429 279457
rect 120371 278969 120429 278981
rect 120829 279457 120887 279469
rect 120829 278981 120841 279457
rect 120875 278981 120887 279457
rect 120829 278969 120887 278981
rect 121071 279457 121129 279469
rect 121071 278981 121083 279457
rect 121117 278981 121129 279457
rect 121071 278969 121129 278981
rect 121529 279457 121587 279469
rect 121529 278981 121541 279457
rect 121575 278981 121587 279457
rect 121529 278969 121587 278981
rect 120371 278673 120429 278685
rect 120371 278197 120383 278673
rect 120417 278197 120429 278673
rect 120371 278185 120429 278197
rect 120829 278673 120887 278685
rect 120829 278197 120841 278673
rect 120875 278197 120887 278673
rect 120829 278185 120887 278197
rect 121071 278673 121129 278685
rect 121071 278197 121083 278673
rect 121117 278197 121129 278673
rect 121071 278185 121129 278197
rect 121529 278673 121587 278685
rect 121529 278197 121541 278673
rect 121575 278197 121587 278673
rect 121529 278185 121587 278197
rect 120371 277889 120429 277901
rect 120371 277413 120383 277889
rect 120417 277413 120429 277889
rect 120371 277401 120429 277413
rect 120829 277889 120887 277901
rect 120829 277413 120841 277889
rect 120875 277413 120887 277889
rect 120829 277401 120887 277413
rect 121071 277889 121129 277901
rect 121071 277413 121083 277889
rect 121117 277413 121129 277889
rect 121071 277401 121129 277413
rect 121529 277889 121587 277901
rect 121529 277413 121541 277889
rect 121575 277413 121587 277889
rect 121529 277401 121587 277413
rect 120371 277105 120429 277117
rect 120371 276629 120383 277105
rect 120417 276629 120429 277105
rect 120371 276617 120429 276629
rect 120829 277105 120887 277117
rect 120829 276629 120841 277105
rect 120875 276629 120887 277105
rect 120829 276617 120887 276629
rect 121071 277105 121129 277117
rect 121071 276629 121083 277105
rect 121117 276629 121129 277105
rect 121071 276617 121129 276629
rect 121529 277105 121587 277117
rect 121529 276629 121541 277105
rect 121575 276629 121587 277105
rect 121529 276617 121587 276629
rect 120371 276321 120429 276333
rect 120371 275845 120383 276321
rect 120417 275845 120429 276321
rect 120371 275833 120429 275845
rect 120829 276321 120887 276333
rect 120829 275845 120841 276321
rect 120875 275845 120887 276321
rect 120829 275833 120887 275845
rect 121071 276321 121129 276333
rect 121071 275845 121083 276321
rect 121117 275845 121129 276321
rect 121071 275833 121129 275845
rect 121529 276321 121587 276333
rect 121529 275845 121541 276321
rect 121575 275845 121587 276321
rect 121529 275833 121587 275845
rect 120371 275537 120429 275549
rect 120371 275061 120383 275537
rect 120417 275061 120429 275537
rect 120371 275049 120429 275061
rect 120829 275537 120887 275549
rect 120829 275061 120841 275537
rect 120875 275061 120887 275537
rect 120829 275049 120887 275061
rect 121071 275537 121129 275549
rect 121071 275061 121083 275537
rect 121117 275061 121129 275537
rect 121071 275049 121129 275061
rect 121529 275537 121587 275549
rect 121529 275061 121541 275537
rect 121575 275061 121587 275537
rect 121529 275049 121587 275061
rect 120371 274753 120429 274765
rect 120371 274277 120383 274753
rect 120417 274277 120429 274753
rect 120371 274265 120429 274277
rect 120829 274753 120887 274765
rect 120829 274277 120841 274753
rect 120875 274277 120887 274753
rect 120829 274265 120887 274277
rect 121071 274753 121129 274765
rect 121071 274277 121083 274753
rect 121117 274277 121129 274753
rect 121071 274265 121129 274277
rect 121529 274753 121587 274765
rect 121529 274277 121541 274753
rect 121575 274277 121587 274753
rect 121529 274265 121587 274277
rect 120371 273969 120429 273981
rect 120371 273493 120383 273969
rect 120417 273493 120429 273969
rect 120371 273481 120429 273493
rect 120829 273969 120887 273981
rect 120829 273493 120841 273969
rect 120875 273493 120887 273969
rect 120829 273481 120887 273493
rect 121071 273969 121129 273981
rect 121071 273493 121083 273969
rect 121117 273493 121129 273969
rect 121071 273481 121129 273493
rect 121529 273969 121587 273981
rect 121529 273493 121541 273969
rect 121575 273493 121587 273969
rect 121529 273481 121587 273493
rect 120371 273185 120429 273197
rect 120371 272709 120383 273185
rect 120417 272709 120429 273185
rect 120371 272697 120429 272709
rect 120829 273185 120887 273197
rect 120829 272709 120841 273185
rect 120875 272709 120887 273185
rect 120829 272697 120887 272709
rect 121071 273185 121129 273197
rect 121071 272709 121083 273185
rect 121117 272709 121129 273185
rect 121071 272697 121129 272709
rect 121529 273185 121587 273197
rect 121529 272709 121541 273185
rect 121575 272709 121587 273185
rect 121529 272697 121587 272709
rect 120371 272401 120429 272413
rect 120371 271925 120383 272401
rect 120417 271925 120429 272401
rect 120371 271913 120429 271925
rect 120829 272401 120887 272413
rect 120829 271925 120841 272401
rect 120875 271925 120887 272401
rect 120829 271913 120887 271925
rect 121071 272401 121129 272413
rect 121071 271925 121083 272401
rect 121117 271925 121129 272401
rect 121071 271913 121129 271925
rect 121529 272401 121587 272413
rect 121529 271925 121541 272401
rect 121575 271925 121587 272401
rect 121529 271913 121587 271925
rect 120371 271617 120429 271629
rect 120371 271141 120383 271617
rect 120417 271141 120429 271617
rect 120371 271129 120429 271141
rect 120829 271617 120887 271629
rect 120829 271141 120841 271617
rect 120875 271141 120887 271617
rect 120829 271129 120887 271141
rect 121071 271617 121129 271629
rect 121071 271141 121083 271617
rect 121117 271141 121129 271617
rect 121071 271129 121129 271141
rect 121529 271617 121587 271629
rect 121529 271141 121541 271617
rect 121575 271141 121587 271617
rect 121529 271129 121587 271141
rect 120371 270833 120429 270845
rect 120371 270357 120383 270833
rect 120417 270357 120429 270833
rect 120371 270345 120429 270357
rect 120829 270833 120887 270845
rect 120829 270357 120841 270833
rect 120875 270357 120887 270833
rect 120829 270345 120887 270357
rect 121071 270833 121129 270845
rect 121071 270357 121083 270833
rect 121117 270357 121129 270833
rect 121071 270345 121129 270357
rect 121529 270833 121587 270845
rect 121529 270357 121541 270833
rect 121575 270357 121587 270833
rect 121529 270345 121587 270357
rect 120371 270049 120429 270061
rect 120371 269573 120383 270049
rect 120417 269573 120429 270049
rect 120371 269561 120429 269573
rect 120829 270049 120887 270061
rect 120829 269573 120841 270049
rect 120875 269573 120887 270049
rect 120829 269561 120887 269573
rect 121071 270049 121129 270061
rect 121071 269573 121083 270049
rect 121117 269573 121129 270049
rect 121071 269561 121129 269573
rect 121529 270049 121587 270061
rect 121529 269573 121541 270049
rect 121575 269573 121587 270049
rect 121529 269561 121587 269573
rect 120371 269265 120429 269277
rect 120371 269189 120383 269265
rect 120417 269189 120429 269265
rect 120371 269177 120429 269189
rect 120829 269265 120887 269277
rect 120829 269189 120841 269265
rect 120875 269189 120887 269265
rect 120829 269177 120887 269189
rect 121071 269265 121129 269277
rect 121071 269189 121083 269265
rect 121117 269189 121129 269265
rect 121071 269177 121129 269189
rect 121529 269265 121587 269277
rect 121529 269189 121541 269265
rect 121575 269189 121587 269265
rect 121529 269177 121587 269189
rect 122298 280411 122356 280423
rect 122298 279935 122310 280411
rect 122344 279935 122356 280411
rect 122298 279923 122356 279935
rect 122756 280411 122814 280423
rect 122756 279935 122768 280411
rect 122802 279935 122814 280411
rect 122756 279923 122814 279935
rect 122998 280411 123056 280423
rect 122998 279935 123010 280411
rect 123044 279935 123056 280411
rect 122998 279923 123056 279935
rect 123456 280411 123514 280423
rect 123456 279935 123468 280411
rect 123502 279935 123514 280411
rect 123456 279923 123514 279935
rect 122298 279627 122356 279639
rect 122298 279151 122310 279627
rect 122344 279151 122356 279627
rect 122298 279139 122356 279151
rect 122756 279627 122814 279639
rect 122756 279151 122768 279627
rect 122802 279151 122814 279627
rect 122756 279139 122814 279151
rect 122998 279627 123056 279639
rect 122998 279151 123010 279627
rect 123044 279151 123056 279627
rect 122998 279139 123056 279151
rect 123456 279627 123514 279639
rect 123456 279151 123468 279627
rect 123502 279151 123514 279627
rect 123456 279139 123514 279151
rect 122356 278254 122414 278266
rect 122356 277804 122368 278254
rect 122402 277804 122414 278254
rect 122356 277792 122414 277804
rect 123290 278254 123348 278266
rect 123290 277804 123302 278254
rect 123336 277804 123348 278254
rect 123290 277792 123348 277804
rect 123598 278068 123656 278080
rect 122358 277488 122416 277500
rect 122358 277412 122370 277488
rect 122404 277412 122416 277488
rect 122358 277400 122416 277412
rect 123216 277488 123274 277500
rect 123216 277412 123228 277488
rect 123262 277412 123274 277488
rect 123216 277400 123274 277412
rect 123598 277406 123610 278068
rect 123644 277406 123656 278068
rect 123598 277394 123656 277406
rect 124210 278068 124268 278080
rect 124210 277406 124222 278068
rect 124256 277406 124268 278068
rect 124210 277394 124268 277406
rect 122380 276656 122438 276668
rect 122380 276504 122392 276656
rect 122426 276504 122438 276656
rect 122380 276492 122438 276504
rect 123832 276656 123890 276668
rect 123832 276504 123844 276656
rect 123878 276504 123890 276656
rect 123832 276492 123890 276504
rect 122466 275857 122866 275869
rect 122466 275823 122478 275857
rect 122854 275823 122866 275857
rect 122466 275811 122866 275823
rect 123102 275857 123502 275869
rect 123102 275823 123114 275857
rect 123490 275823 123502 275857
rect 123102 275811 123502 275823
rect 123738 275857 124138 275869
rect 123738 275823 123750 275857
rect 124126 275823 124138 275857
rect 123738 275811 124138 275823
rect 124374 275857 124774 275869
rect 124374 275823 124386 275857
rect 124762 275823 124774 275857
rect 124374 275811 124774 275823
rect 122466 275699 122866 275711
rect 122466 275665 122478 275699
rect 122854 275665 122866 275699
rect 122466 275653 122866 275665
rect 123102 275699 123502 275711
rect 123102 275665 123114 275699
rect 123490 275665 123502 275699
rect 123102 275653 123502 275665
rect 123738 275699 124138 275711
rect 123738 275665 123750 275699
rect 124126 275665 124138 275699
rect 123738 275653 124138 275665
rect 124374 275699 124774 275711
rect 124374 275665 124386 275699
rect 124762 275665 124774 275699
rect 124374 275653 124774 275665
rect 122067 272801 122125 272813
rect 122067 272725 122079 272801
rect 122113 272725 122125 272801
rect 122067 272713 122125 272725
rect 122525 272801 122583 272813
rect 122525 272725 122537 272801
rect 122571 272725 122583 272801
rect 122525 272713 122583 272725
rect 122767 272801 122825 272813
rect 122767 272725 122779 272801
rect 122813 272725 122825 272801
rect 122767 272713 122825 272725
rect 123225 272801 123283 272813
rect 123225 272725 123237 272801
rect 123271 272725 123283 272801
rect 123225 272713 123283 272725
rect 122067 272417 122125 272429
rect 122067 271941 122079 272417
rect 122113 271941 122125 272417
rect 122067 271929 122125 271941
rect 122525 272417 122583 272429
rect 122525 271941 122537 272417
rect 122571 271941 122583 272417
rect 122525 271929 122583 271941
rect 122767 272417 122825 272429
rect 122767 271941 122779 272417
rect 122813 271941 122825 272417
rect 122767 271929 122825 271941
rect 123225 272417 123283 272429
rect 123225 271941 123237 272417
rect 123271 271941 123283 272417
rect 123225 271929 123283 271941
rect 122067 271633 122125 271645
rect 122067 271157 122079 271633
rect 122113 271157 122125 271633
rect 122067 271145 122125 271157
rect 122525 271633 122583 271645
rect 122525 271157 122537 271633
rect 122571 271157 122583 271633
rect 122525 271145 122583 271157
rect 122767 271633 122825 271645
rect 122767 271157 122779 271633
rect 122813 271157 122825 271633
rect 122767 271145 122825 271157
rect 123225 271633 123283 271645
rect 123225 271157 123237 271633
rect 123271 271157 123283 271633
rect 123225 271145 123283 271157
rect 122067 270849 122125 270861
rect 122067 270373 122079 270849
rect 122113 270373 122125 270849
rect 122067 270361 122125 270373
rect 122525 270849 122583 270861
rect 122525 270373 122537 270849
rect 122571 270373 122583 270849
rect 122525 270361 122583 270373
rect 122767 270849 122825 270861
rect 122767 270373 122779 270849
rect 122813 270373 122825 270849
rect 122767 270361 122825 270373
rect 123225 270849 123283 270861
rect 123225 270373 123237 270849
rect 123271 270373 123283 270849
rect 123225 270361 123283 270373
rect 122067 270065 122125 270077
rect 122067 269589 122079 270065
rect 122113 269589 122125 270065
rect 122067 269577 122125 269589
rect 122525 270065 122583 270077
rect 122525 269589 122537 270065
rect 122571 269589 122583 270065
rect 122525 269577 122583 269589
rect 122767 270065 122825 270077
rect 122767 269589 122779 270065
rect 122813 269589 122825 270065
rect 122767 269577 122825 269589
rect 123225 270065 123283 270077
rect 123225 269589 123237 270065
rect 123271 269589 123283 270065
rect 123225 269577 123283 269589
rect 122067 269281 122125 269293
rect 122067 269205 122079 269281
rect 122113 269205 122125 269281
rect 122067 269193 122125 269205
rect 122525 269281 122583 269293
rect 122525 269205 122537 269281
rect 122571 269205 122583 269281
rect 122525 269193 122583 269205
rect 122767 269281 122825 269293
rect 122767 269205 122779 269281
rect 122813 269205 122825 269281
rect 122767 269193 122825 269205
rect 123225 269281 123283 269293
rect 123225 269205 123237 269281
rect 123271 269205 123283 269281
rect 123225 269193 123283 269205
<< ndiffc >>
rect 106311 279805 106345 280801
rect 106501 279805 106535 280801
rect 106711 279805 106745 280801
rect 106901 279805 106935 280801
rect 107111 279805 107145 280801
rect 107301 279805 107335 280801
rect 107511 279805 107545 280801
rect 107701 279805 107735 280801
rect 107911 279805 107945 280801
rect 108101 279805 108135 280801
rect 108311 279805 108345 280801
rect 108501 279805 108535 280801
rect 108711 279805 108745 280801
rect 108901 279805 108935 280801
rect 109111 279805 109145 280801
rect 109301 279805 109335 280801
rect 109511 279805 109545 280801
rect 109701 279805 109735 280801
rect 109911 279805 109945 280801
rect 110101 279805 110135 280801
rect 109731 277985 109765 278999
rect 110075 277985 110109 278999
rect 109731 276729 109765 277743
rect 110075 276729 110109 277743
rect 106935 271819 106969 271959
rect 107203 271819 107237 271959
rect 107413 271747 107447 272067
rect 108091 271747 108125 272067
rect 107185 271501 108361 271535
rect 107185 271265 108361 271299
rect 107185 271131 108361 271165
rect 107185 270895 108361 270929
rect 111536 280832 112612 280866
rect 112982 280840 114058 280874
rect 111536 280614 112612 280648
rect 112982 280582 114058 280616
rect 111536 280472 112612 280506
rect 112982 280416 114058 280450
rect 111536 280254 112612 280288
rect 112982 280158 114058 280192
rect 111536 280112 112612 280146
rect 113012 280014 114088 280048
rect 111536 279894 112612 279928
rect 113012 279876 114088 279910
rect 111536 279752 112612 279786
rect 113012 279716 114088 279750
rect 111536 279534 112612 279568
rect 113012 279578 114088 279612
rect 116147 280840 117223 280874
rect 117593 280832 118669 280866
rect 116147 280582 117223 280616
rect 117593 280614 118669 280648
rect 117593 280472 118669 280506
rect 116147 280416 117223 280450
rect 117593 280254 118669 280288
rect 116147 280158 117223 280192
rect 117593 280112 118669 280146
rect 116117 280014 117193 280048
rect 116117 279876 117193 279910
rect 117593 279894 118669 279928
rect 116117 279716 117193 279750
rect 117593 279752 118669 279786
rect 116117 279578 117193 279612
rect 117593 279534 118669 279568
rect 111536 279166 112612 279200
rect 112982 279174 114058 279208
rect 111536 278948 112612 278982
rect 112982 278916 114058 278950
rect 111536 278806 112612 278840
rect 112982 278750 114058 278784
rect 111536 278588 112612 278622
rect 112982 278492 114058 278526
rect 111536 278446 112612 278480
rect 113012 278348 114088 278382
rect 111536 278228 112612 278262
rect 113012 278210 114088 278244
rect 111536 278086 112612 278120
rect 113012 278050 114088 278084
rect 111536 277868 112612 277902
rect 113012 277912 114088 277946
rect 116147 279174 117223 279208
rect 117593 279166 118669 279200
rect 116147 278916 117223 278950
rect 117593 278948 118669 278982
rect 117593 278806 118669 278840
rect 116147 278750 117223 278784
rect 117593 278588 118669 278622
rect 116147 278492 117223 278526
rect 117593 278446 118669 278480
rect 116117 278348 117193 278382
rect 116117 278210 117193 278244
rect 117593 278228 118669 278262
rect 116117 278050 117193 278084
rect 117593 278086 118669 278120
rect 116117 277912 117193 277946
rect 117593 277868 118669 277902
rect 111536 277500 112612 277534
rect 112982 277508 114058 277542
rect 111536 277282 112612 277316
rect 112982 277250 114058 277284
rect 111536 277140 112612 277174
rect 112982 277084 114058 277118
rect 111536 276922 112612 276956
rect 112982 276826 114058 276860
rect 111536 276780 112612 276814
rect 113012 276682 114088 276716
rect 111536 276562 112612 276596
rect 113012 276544 114088 276578
rect 111536 276420 112612 276454
rect 113012 276384 114088 276418
rect 111536 276202 112612 276236
rect 113012 276246 114088 276280
rect 116147 277508 117223 277542
rect 117593 277500 118669 277534
rect 116147 277250 117223 277284
rect 117593 277282 118669 277316
rect 117593 277140 118669 277174
rect 116147 277084 117223 277118
rect 117593 276922 118669 276956
rect 116147 276826 117223 276860
rect 117593 276780 118669 276814
rect 116117 276682 117193 276716
rect 116117 276544 117193 276578
rect 117593 276562 118669 276596
rect 116117 276384 117193 276418
rect 117593 276420 118669 276454
rect 116117 276246 117193 276280
rect 117593 276202 118669 276236
rect 111536 275834 112612 275868
rect 112982 275842 114058 275876
rect 111536 275616 112612 275650
rect 112982 275584 114058 275618
rect 111536 275474 112612 275508
rect 112982 275418 114058 275452
rect 111536 275256 112612 275290
rect 112982 275160 114058 275194
rect 111536 275114 112612 275148
rect 113012 275016 114088 275050
rect 111536 274896 112612 274930
rect 113012 274878 114088 274912
rect 111536 274754 112612 274788
rect 113012 274718 114088 274752
rect 111536 274536 112612 274570
rect 113012 274580 114088 274614
rect 116147 275842 117223 275876
rect 117593 275834 118669 275868
rect 116147 275584 117223 275618
rect 117593 275616 118669 275650
rect 117593 275474 118669 275508
rect 116147 275418 117223 275452
rect 117593 275256 118669 275290
rect 116147 275160 117223 275194
rect 117593 275114 118669 275148
rect 116117 275016 117193 275050
rect 116117 274878 117193 274912
rect 117593 274896 118669 274930
rect 116117 274718 117193 274752
rect 117593 274754 118669 274788
rect 116117 274580 117193 274614
rect 117593 274536 118669 274570
rect 111536 274168 112612 274202
rect 112982 274176 114058 274210
rect 111536 273950 112612 273984
rect 112982 273918 114058 273952
rect 111536 273808 112612 273842
rect 112982 273752 114058 273786
rect 111536 273590 112612 273624
rect 112982 273494 114058 273528
rect 111536 273448 112612 273482
rect 113012 273350 114088 273384
rect 111536 273230 112612 273264
rect 113012 273212 114088 273246
rect 111536 273088 112612 273122
rect 113012 273052 114088 273086
rect 111536 272870 112612 272904
rect 113012 272914 114088 272948
rect 116147 274176 117223 274210
rect 117593 274168 118669 274202
rect 116147 273918 117223 273952
rect 117593 273950 118669 273984
rect 117593 273808 118669 273842
rect 116147 273752 117223 273786
rect 117593 273590 118669 273624
rect 116147 273494 117223 273528
rect 117593 273448 118669 273482
rect 116117 273350 117193 273384
rect 116117 273212 117193 273246
rect 117593 273230 118669 273264
rect 116117 273052 117193 273086
rect 117593 273088 118669 273122
rect 116117 272914 117193 272948
rect 117593 272870 118669 272904
rect 115835 270836 115869 271912
rect 116053 270836 116087 271912
rect 116235 270836 116269 271912
rect 116453 270836 116487 271912
rect 116635 270836 116669 271912
rect 116853 270836 116887 271912
rect 117035 270836 117069 271912
rect 117253 270836 117287 271912
rect 117435 270836 117469 271912
rect 117653 270836 117687 271912
rect 117835 270836 117869 271912
rect 118053 270836 118087 271912
rect 118235 270836 118269 271912
rect 118453 270836 118487 271912
rect 118635 270836 118669 271912
rect 118853 270836 118887 271912
rect 112514 269136 112548 270212
rect 112732 269136 112766 270212
rect 112914 269136 112948 270212
rect 113132 269136 113166 270212
rect 113314 269136 113348 270212
rect 113532 269136 113566 270212
rect 113714 269136 113748 270212
rect 113932 269136 113966 270212
rect 114114 269136 114148 270212
rect 114332 269136 114366 270212
rect 114514 269136 114548 270212
rect 114732 269136 114766 270212
rect 114914 269136 114948 270212
rect 115132 269136 115166 270212
rect 115314 269136 115348 270212
rect 115532 269136 115566 270212
rect 115714 269136 115748 270212
rect 115932 269136 115966 270212
rect 116114 269136 116148 270212
rect 116332 269136 116366 270212
rect 116514 269136 116548 270212
rect 116732 269136 116766 270212
rect 116914 269136 116948 270212
rect 117132 269136 117166 270212
rect 117314 269136 117348 270212
rect 117532 269136 117566 270212
rect 117714 269136 117748 270212
rect 117932 269136 117966 270212
rect 118114 269136 118148 270212
rect 118332 269136 118366 270212
rect 118514 269136 118548 270212
rect 118732 269136 118766 270212
rect 122906 274674 122940 274850
rect 123964 274674 123998 274850
rect 122231 273790 122265 274266
rect 122489 273790 122523 274266
rect 122647 273790 122681 274266
rect 122905 273790 122939 274266
rect 123063 273790 123097 274266
rect 123321 273790 123355 274266
rect 123479 273790 123513 274266
rect 123737 273790 123771 274266
rect 123895 273790 123929 274266
rect 124153 273790 124187 274266
rect 124311 273790 124345 274266
rect 124569 273790 124603 274266
rect 124204 272532 124680 272566
rect 124204 272274 124680 272308
rect 124204 272116 124680 272150
rect 124204 271858 124680 271892
rect 124204 271700 124680 271734
rect 124204 271442 124680 271476
rect 124204 271284 124680 271318
rect 124204 271026 124680 271060
rect 124204 270868 124680 270902
rect 124204 270610 124680 270644
rect 124204 270452 124680 270486
rect 124204 270194 124680 270228
rect 124204 270036 124680 270070
rect 124204 269778 124680 269812
rect 124204 269620 124680 269654
rect 124204 269362 124680 269396
<< pdiffc >>
rect 106380 279023 107570 279057
rect 106380 278711 107570 278745
rect 106380 278423 107570 278457
rect 106380 278111 107570 278145
rect 106503 277176 107513 277210
rect 106503 277044 107513 277078
rect 106963 275725 107117 275759
rect 107463 275725 107617 275759
rect 107963 275725 108117 275759
rect 108463 275725 108617 275759
rect 108963 275725 109117 275759
rect 109463 275725 109617 275759
rect 106963 274889 107117 274923
rect 107463 274889 107617 274923
rect 107963 274889 108117 274923
rect 108463 274889 108617 274923
rect 108963 274889 109117 274923
rect 109463 274889 109617 274923
rect 109394 270718 109428 272414
rect 109522 270718 109556 272414
rect 114669 280815 114845 280849
rect 114669 280357 114845 280391
rect 114669 280129 114845 280163
rect 114669 279911 114845 279945
rect 114669 279721 114845 279755
rect 114669 279503 114845 279537
rect 115360 280815 115536 280849
rect 115360 280357 115536 280391
rect 115360 280129 115536 280163
rect 115360 279911 115536 279945
rect 115360 279721 115536 279755
rect 115360 279503 115536 279537
rect 114669 279149 114845 279183
rect 114669 278691 114845 278725
rect 114669 278463 114845 278497
rect 114669 278245 114845 278279
rect 114669 278055 114845 278089
rect 114669 277837 114845 277871
rect 115360 279149 115536 279183
rect 115360 278691 115536 278725
rect 115360 278463 115536 278497
rect 115360 278245 115536 278279
rect 115360 278055 115536 278089
rect 115360 277837 115536 277871
rect 114669 277483 114845 277517
rect 114669 277025 114845 277059
rect 114669 276797 114845 276831
rect 114669 276579 114845 276613
rect 114669 276389 114845 276423
rect 114669 276171 114845 276205
rect 115360 277483 115536 277517
rect 115360 277025 115536 277059
rect 115360 276797 115536 276831
rect 115360 276579 115536 276613
rect 115360 276389 115536 276423
rect 115360 276171 115536 276205
rect 114669 275817 114845 275851
rect 114669 275359 114845 275393
rect 114669 275131 114845 275165
rect 114669 274913 114845 274947
rect 114669 274723 114845 274757
rect 114669 274505 114845 274539
rect 115360 275817 115536 275851
rect 115360 275359 115536 275393
rect 115360 275131 115536 275165
rect 115360 274913 115536 274947
rect 115360 274723 115536 274757
rect 115360 274505 115536 274539
rect 114669 274151 114845 274185
rect 114669 273693 114845 273727
rect 114669 273465 114845 273499
rect 114669 273247 114845 273281
rect 114669 273057 114845 273091
rect 114669 272839 114845 272873
rect 115360 274151 115536 274185
rect 115360 273693 115536 273727
rect 115360 273465 115536 273499
rect 115360 273247 115536 273281
rect 115360 273057 115536 273091
rect 115360 272839 115536 272873
rect 112532 271118 112566 271294
rect 112750 271118 112784 271294
rect 112932 271118 112966 271294
rect 113150 271118 113184 271294
rect 113332 271118 113366 271294
rect 113550 271118 113584 271294
rect 113732 271118 113766 271294
rect 113950 271118 113984 271294
rect 114591 271089 114625 271265
rect 114809 271089 114843 271265
rect 114991 271089 115025 271265
rect 115209 271089 115243 271265
rect 120383 280549 120417 280625
rect 120841 280549 120875 280625
rect 121083 280549 121117 280625
rect 121541 280549 121575 280625
rect 120383 279765 120417 280241
rect 120841 279765 120875 280241
rect 121083 279765 121117 280241
rect 121541 279765 121575 280241
rect 120383 278981 120417 279457
rect 120841 278981 120875 279457
rect 121083 278981 121117 279457
rect 121541 278981 121575 279457
rect 120383 278197 120417 278673
rect 120841 278197 120875 278673
rect 121083 278197 121117 278673
rect 121541 278197 121575 278673
rect 120383 277413 120417 277889
rect 120841 277413 120875 277889
rect 121083 277413 121117 277889
rect 121541 277413 121575 277889
rect 120383 276629 120417 277105
rect 120841 276629 120875 277105
rect 121083 276629 121117 277105
rect 121541 276629 121575 277105
rect 120383 275845 120417 276321
rect 120841 275845 120875 276321
rect 121083 275845 121117 276321
rect 121541 275845 121575 276321
rect 120383 275061 120417 275537
rect 120841 275061 120875 275537
rect 121083 275061 121117 275537
rect 121541 275061 121575 275537
rect 120383 274277 120417 274753
rect 120841 274277 120875 274753
rect 121083 274277 121117 274753
rect 121541 274277 121575 274753
rect 120383 273493 120417 273969
rect 120841 273493 120875 273969
rect 121083 273493 121117 273969
rect 121541 273493 121575 273969
rect 120383 272709 120417 273185
rect 120841 272709 120875 273185
rect 121083 272709 121117 273185
rect 121541 272709 121575 273185
rect 120383 271925 120417 272401
rect 120841 271925 120875 272401
rect 121083 271925 121117 272401
rect 121541 271925 121575 272401
rect 120383 271141 120417 271617
rect 120841 271141 120875 271617
rect 121083 271141 121117 271617
rect 121541 271141 121575 271617
rect 120383 270357 120417 270833
rect 120841 270357 120875 270833
rect 121083 270357 121117 270833
rect 121541 270357 121575 270833
rect 120383 269573 120417 270049
rect 120841 269573 120875 270049
rect 121083 269573 121117 270049
rect 121541 269573 121575 270049
rect 120383 269189 120417 269265
rect 120841 269189 120875 269265
rect 121083 269189 121117 269265
rect 121541 269189 121575 269265
rect 122310 279935 122344 280411
rect 122768 279935 122802 280411
rect 123010 279935 123044 280411
rect 123468 279935 123502 280411
rect 122310 279151 122344 279627
rect 122768 279151 122802 279627
rect 123010 279151 123044 279627
rect 123468 279151 123502 279627
rect 122368 277804 122402 278254
rect 123302 277804 123336 278254
rect 122370 277412 122404 277488
rect 123228 277412 123262 277488
rect 123610 277406 123644 278068
rect 124222 277406 124256 278068
rect 122392 276504 122426 276656
rect 123844 276504 123878 276656
rect 122478 275823 122854 275857
rect 123114 275823 123490 275857
rect 123750 275823 124126 275857
rect 124386 275823 124762 275857
rect 122478 275665 122854 275699
rect 123114 275665 123490 275699
rect 123750 275665 124126 275699
rect 124386 275665 124762 275699
rect 122079 272725 122113 272801
rect 122537 272725 122571 272801
rect 122779 272725 122813 272801
rect 123237 272725 123271 272801
rect 122079 271941 122113 272417
rect 122537 271941 122571 272417
rect 122779 271941 122813 272417
rect 123237 271941 123271 272417
rect 122079 271157 122113 271633
rect 122537 271157 122571 271633
rect 122779 271157 122813 271633
rect 123237 271157 123271 271633
rect 122079 270373 122113 270849
rect 122537 270373 122571 270849
rect 122779 270373 122813 270849
rect 123237 270373 123271 270849
rect 122079 269589 122113 270065
rect 122537 269589 122571 270065
rect 122779 269589 122813 270065
rect 123237 269589 123271 270065
rect 122079 269205 122113 269281
rect 122537 269205 122571 269281
rect 122779 269205 122813 269281
rect 123237 269205 123271 269281
<< psubdiff >>
rect 111046 281107 111234 281179
rect 105974 281045 106147 281065
rect 105974 281041 106170 281045
rect 106060 280961 106170 281041
rect 110228 280961 110313 281045
rect 106060 280880 106207 280961
rect 106060 279716 106125 280880
rect 110231 280862 110313 280961
rect 106060 279625 106207 279716
rect 110231 279625 110313 279698
rect 106060 279541 106170 279625
rect 110228 279541 110313 279625
rect 110053 279185 110187 279541
rect 109617 279151 109713 279185
rect 110127 279151 110223 279185
rect 109617 279089 109651 279151
rect 110189 279089 110223 279151
rect 109617 276577 109651 276639
rect 110189 276577 110223 276639
rect 109617 276543 109713 276577
rect 110127 276548 110223 276577
rect 110127 276543 110224 276548
rect 110145 276056 110224 276543
rect 105974 274619 106060 274635
rect 110145 274619 110224 274669
rect 105974 274527 106114 274619
rect 110167 274527 110224 274619
rect 106281 272918 106580 272951
rect 106459 272794 106580 272918
rect 109977 272918 110259 272951
rect 109977 272794 110081 272918
rect 106459 272786 110081 272794
rect 106715 272339 106843 272367
rect 106789 272299 106843 272339
rect 106887 272299 106963 272367
rect 108657 272339 108803 272367
rect 108657 272299 108729 272339
rect 106789 270773 106869 270801
rect 106715 270733 106869 270773
rect 108683 270773 108729 270801
rect 108683 270733 108803 270773
rect 106459 270193 106570 270334
rect 106281 270177 106570 270193
rect 109967 270193 110081 270334
rect 111200 281099 111234 281107
rect 118876 281107 119159 281179
rect 118876 281099 119005 281107
rect 114235 280884 114353 280908
rect 114235 280742 114353 280766
rect 111200 279335 111328 279425
rect 114242 279335 114266 279425
rect 115852 280884 115970 280908
rect 115852 280742 115970 280766
rect 115939 279335 115963 279425
rect 118877 279335 119005 279425
rect 114235 279218 114353 279242
rect 114235 279076 114353 279100
rect 111200 277669 111328 277759
rect 114242 277669 114266 277759
rect 115852 279218 115970 279242
rect 115852 279076 115970 279100
rect 115939 277669 115963 277759
rect 118877 277669 119005 277759
rect 114235 277552 114353 277576
rect 114235 277410 114353 277434
rect 111200 276003 111328 276093
rect 114242 276003 114266 276093
rect 115852 277552 115970 277576
rect 115852 277410 115970 277434
rect 115939 276003 115963 276093
rect 118877 276003 119005 276093
rect 114235 275886 114353 275910
rect 114235 275744 114353 275768
rect 111200 274337 111328 274427
rect 114242 274337 114266 274427
rect 115852 275886 115970 275910
rect 115852 275744 115970 275768
rect 115939 274337 115963 274427
rect 118877 274337 119005 274427
rect 114235 274220 114353 274244
rect 114235 274078 114353 274102
rect 114143 272761 114266 272766
rect 111200 272699 111328 272761
rect 111046 272671 111328 272699
rect 114242 272671 114266 272761
rect 115852 274220 115970 274244
rect 115852 274078 115970 274102
rect 115939 272761 116062 272766
rect 114143 272551 114266 272671
rect 115939 272671 115963 272761
rect 118877 272699 119005 272761
rect 118877 272671 119159 272699
rect 119938 281067 120227 281165
rect 115939 272551 116062 272671
rect 114143 272460 116062 272551
rect 109967 270177 110259 270193
rect 106281 270169 110259 270177
rect 111939 272249 112069 272273
rect 119021 272249 119151 272273
rect 112069 272125 112167 272249
rect 118956 272125 119021 272249
rect 112069 268702 112160 268826
rect 118949 268702 119021 268826
rect 111939 268651 112069 268675
rect 120104 281012 120227 281067
rect 125148 281012 125172 281165
rect 125047 280856 125171 281012
rect 122027 278619 122144 278643
rect 122144 276097 122500 276212
rect 124297 276097 124321 276212
rect 122027 275507 122144 275531
rect 122792 275002 122888 275036
rect 124016 275002 124112 275036
rect 122792 274940 122826 275002
rect 124078 274940 124112 275002
rect 122792 274562 122826 274584
rect 124078 274582 124112 274584
rect 122060 274486 122084 274562
rect 122714 274522 122826 274562
rect 124078 274522 124218 274582
rect 122714 274488 122888 274522
rect 124016 274488 124218 274522
rect 124824 274488 124848 274582
rect 122714 274486 122807 274488
rect 122060 274384 122150 274486
rect 122062 274296 122150 274384
rect 124726 274312 124814 274488
rect 122062 273618 122150 273621
rect 124726 273618 124814 273637
rect 122062 273545 122217 273618
rect 124615 273545 124814 273618
rect 123978 272689 124051 272777
rect 124726 272717 124880 272777
rect 124726 272689 124811 272717
rect 123978 272598 124029 272689
rect 123978 269281 124029 269356
rect 124811 269281 124880 269291
rect 123978 269193 124035 269281
rect 124710 269193 124880 269281
rect 125047 268861 125171 268990
rect 120104 268778 120254 268861
rect 119938 268708 120254 268778
rect 125175 268708 125199 268861
rect 119021 268651 119151 268675
<< nsubdiff >>
rect 106169 279188 106229 279222
rect 107708 279188 107768 279222
rect 106169 279162 106203 279188
rect 107734 279162 107768 279188
rect 106169 277984 106203 278010
rect 107734 277984 107768 278010
rect 106169 277950 106229 277984
rect 107708 277950 107768 277984
rect 106308 277290 106404 277324
rect 107612 277290 107708 277324
rect 106308 277228 106342 277290
rect 107674 277228 107708 277290
rect 106308 276964 106342 277026
rect 107674 276964 107708 277026
rect 106308 276930 106404 276964
rect 107612 276930 107708 276964
rect 106706 275900 106766 275934
rect 109787 275900 109847 275934
rect 106706 275874 106740 275900
rect 109813 275874 109847 275900
rect 106706 274747 106740 274773
rect 109813 274747 109847 274773
rect 106706 274713 106766 274747
rect 109787 274713 109847 274747
rect 109088 272568 109148 272602
rect 109801 272568 109861 272602
rect 109088 272542 109122 272568
rect 109827 272542 109861 272568
rect 109088 270555 109122 270581
rect 109827 270555 109861 270581
rect 109088 270521 109148 270555
rect 109801 270521 109861 270555
rect 114455 280929 114515 280963
rect 115001 280929 115061 280963
rect 114455 280903 114489 280929
rect 115027 280903 115061 280929
rect 114455 279403 114489 279429
rect 115027 279403 115061 279429
rect 114455 279369 114515 279403
rect 115001 279369 115061 279403
rect 115144 280929 115204 280963
rect 115690 280929 115750 280963
rect 115144 280903 115178 280929
rect 115716 280903 115750 280929
rect 115144 279403 115178 279429
rect 115716 279403 115750 279429
rect 115144 279369 115204 279403
rect 115690 279369 115750 279403
rect 114455 279263 114515 279297
rect 115001 279263 115061 279297
rect 114455 279237 114489 279263
rect 115027 279237 115061 279263
rect 114455 277737 114489 277763
rect 115027 277737 115061 277763
rect 114455 277703 114515 277737
rect 115001 277703 115061 277737
rect 115144 279263 115204 279297
rect 115690 279263 115750 279297
rect 115144 279237 115178 279263
rect 115716 279237 115750 279263
rect 115144 277737 115178 277763
rect 115716 277737 115750 277763
rect 115144 277703 115204 277737
rect 115690 277703 115750 277737
rect 114455 277597 114515 277631
rect 115001 277597 115061 277631
rect 114455 277571 114489 277597
rect 115027 277571 115061 277597
rect 114455 276071 114489 276097
rect 115027 276071 115061 276097
rect 114455 276037 114515 276071
rect 115001 276037 115061 276071
rect 115144 277597 115204 277631
rect 115690 277597 115750 277631
rect 115144 277571 115178 277597
rect 115716 277571 115750 277597
rect 115144 276071 115178 276097
rect 115716 276071 115750 276097
rect 115144 276037 115204 276071
rect 115690 276037 115750 276071
rect 114455 275931 114515 275965
rect 115001 275931 115061 275965
rect 114455 275905 114489 275931
rect 115027 275905 115061 275931
rect 114455 274405 114489 274431
rect 115027 274405 115061 274431
rect 114455 274371 114515 274405
rect 115001 274371 115061 274405
rect 115144 275931 115204 275965
rect 115690 275931 115750 275965
rect 115144 275905 115178 275931
rect 115716 275905 115750 275931
rect 115144 274405 115178 274431
rect 115716 274405 115750 274431
rect 115144 274371 115204 274405
rect 115690 274371 115750 274405
rect 114455 274265 114515 274299
rect 115001 274265 115061 274299
rect 114455 274239 114489 274265
rect 115027 274239 115061 274265
rect 114455 272739 114489 272765
rect 115027 272739 115061 272765
rect 114455 272705 114515 272739
rect 115001 272705 115061 272739
rect 115144 274265 115204 274299
rect 115690 274265 115750 274299
rect 115144 274239 115178 274265
rect 115716 274239 115750 274265
rect 115144 272739 115178 272765
rect 115716 272739 115750 272765
rect 115144 272705 115204 272739
rect 115690 272705 115750 272739
rect 112307 271634 112367 271668
rect 114150 271634 114210 271668
rect 112307 271608 112341 271634
rect 114176 271608 114210 271634
rect 112307 270817 112341 270843
rect 114176 270817 114210 270843
rect 112307 270783 112367 270817
rect 114150 270783 114210 270817
rect 114329 271554 114389 271588
rect 115443 271554 115503 271588
rect 114329 271528 114363 271554
rect 115469 271528 115503 271554
rect 114329 270806 114363 270832
rect 115469 270806 115503 270832
rect 114329 270772 114389 270806
rect 115443 270772 115503 270806
rect 120237 280779 120297 280813
rect 121668 280779 121728 280813
rect 120237 280753 120271 280779
rect 121694 280753 121728 280779
rect 120237 269012 120271 269038
rect 122178 280574 122238 280608
rect 123578 280574 123638 280608
rect 122178 280548 122212 280574
rect 123604 280548 123638 280574
rect 122178 279000 122212 279026
rect 123604 279000 123638 279026
rect 122178 278966 122238 279000
rect 123578 278966 123638 279000
rect 122254 278448 122314 278482
rect 124310 278448 124370 278482
rect 122254 278422 122288 278448
rect 124336 278422 124370 278448
rect 122254 277221 122288 277247
rect 124336 277221 124370 277247
rect 122254 277187 122314 277221
rect 124310 277187 124370 277221
rect 122278 276817 122374 276851
rect 123896 276817 123992 276851
rect 122278 276755 122312 276817
rect 123958 276755 123992 276817
rect 122278 276343 122312 276405
rect 123958 276343 123992 276405
rect 122278 276309 122374 276343
rect 123896 276309 123992 276343
rect 122283 275937 122379 275971
rect 124861 275937 124957 275971
rect 122283 275875 122317 275937
rect 124923 275875 124957 275937
rect 122283 275585 122317 275647
rect 124923 275585 124957 275647
rect 122283 275551 122379 275585
rect 124861 275551 124957 275585
rect 121694 269012 121728 269038
rect 120237 268978 120297 269012
rect 121668 268978 121728 269012
rect 121920 272964 121980 272998
rect 123494 272964 123554 272998
rect 121920 272938 121954 272964
rect 123520 272938 123554 272964
rect 121920 269028 121954 269054
rect 123520 269028 123554 269054
rect 121920 268994 121980 269028
rect 123494 268994 123554 269028
<< psubdiffcont >>
rect 105974 274635 106060 281041
rect 106170 280961 110228 281045
rect 106125 279716 106207 280880
rect 110231 279698 110313 280862
rect 106170 279541 110228 279625
rect 109713 279151 110127 279185
rect 109617 276639 109651 279089
rect 110189 276639 110223 279089
rect 109713 276543 110127 276577
rect 110145 274669 110224 276056
rect 106114 274527 110167 274619
rect 106281 270193 106459 272918
rect 106580 272794 109977 272951
rect 106715 270773 106789 272339
rect 106843 272299 106887 272367
rect 106963 272299 108657 272367
rect 106869 270733 108683 270801
rect 108729 270773 108803 272339
rect 106570 270177 109967 270334
rect 110081 270193 110259 272918
rect 111046 272699 111200 281107
rect 111234 281099 118876 281179
rect 114235 280766 114353 280884
rect 111328 279335 114242 279425
rect 115852 280766 115970 280884
rect 115963 279335 118877 279425
rect 114235 279100 114353 279218
rect 111328 277669 114242 277759
rect 115852 279100 115970 279218
rect 115963 277669 118877 277759
rect 114235 277434 114353 277552
rect 111328 276003 114242 276093
rect 115852 277434 115970 277552
rect 115963 276003 118877 276093
rect 114235 275768 114353 275886
rect 111328 274337 114242 274427
rect 115852 275768 115970 275886
rect 115963 274337 118877 274427
rect 114235 274102 114353 274220
rect 111328 272671 114242 272761
rect 115852 274102 115970 274220
rect 115963 272671 118877 272761
rect 119005 272699 119159 281107
rect 111939 268675 112069 272249
rect 112167 272125 118956 272249
rect 112160 268702 118949 268826
rect 119021 268675 119151 272249
rect 119938 268778 120104 281067
rect 120227 281012 125148 281165
rect 122027 275531 122144 278619
rect 122500 276097 124297 276212
rect 122888 275002 124016 275036
rect 122792 274584 122826 274940
rect 124078 274584 124112 274940
rect 122084 274486 122714 274562
rect 122888 274488 124016 274522
rect 124218 274488 124824 274582
rect 122062 273621 122150 274296
rect 124726 273637 124814 274312
rect 122217 273545 124615 273618
rect 124051 272689 124726 272777
rect 123978 269356 124029 272598
rect 124811 269291 124880 272717
rect 124035 269193 124710 269281
rect 125047 268990 125171 280856
rect 120254 268708 125175 268861
<< nsubdiffcont >>
rect 106229 279188 107708 279222
rect 106169 278010 106203 279162
rect 107734 278010 107768 279162
rect 106229 277950 107708 277984
rect 106404 277290 107612 277324
rect 106308 277026 106342 277228
rect 107674 277026 107708 277228
rect 106404 276930 107612 276964
rect 106766 275900 109787 275934
rect 106706 274773 106740 275874
rect 109813 274773 109847 275874
rect 106766 274713 109787 274747
rect 109148 272568 109801 272602
rect 109088 270581 109122 272542
rect 109827 270581 109861 272542
rect 109148 270521 109801 270555
rect 114515 280929 115001 280963
rect 114455 279429 114489 280903
rect 115027 279429 115061 280903
rect 114515 279369 115001 279403
rect 115204 280929 115690 280963
rect 115144 279429 115178 280903
rect 115716 279429 115750 280903
rect 115204 279369 115690 279403
rect 114515 279263 115001 279297
rect 114455 277763 114489 279237
rect 115027 277763 115061 279237
rect 114515 277703 115001 277737
rect 115204 279263 115690 279297
rect 115144 277763 115178 279237
rect 115716 277763 115750 279237
rect 115204 277703 115690 277737
rect 114515 277597 115001 277631
rect 114455 276097 114489 277571
rect 115027 276097 115061 277571
rect 114515 276037 115001 276071
rect 115204 277597 115690 277631
rect 115144 276097 115178 277571
rect 115716 276097 115750 277571
rect 115204 276037 115690 276071
rect 114515 275931 115001 275965
rect 114455 274431 114489 275905
rect 115027 274431 115061 275905
rect 114515 274371 115001 274405
rect 115204 275931 115690 275965
rect 115144 274431 115178 275905
rect 115716 274431 115750 275905
rect 115204 274371 115690 274405
rect 114515 274265 115001 274299
rect 114455 272765 114489 274239
rect 115027 272765 115061 274239
rect 114515 272705 115001 272739
rect 115204 274265 115690 274299
rect 115144 272765 115178 274239
rect 115716 272765 115750 274239
rect 115204 272705 115690 272739
rect 112367 271634 114150 271668
rect 112307 270843 112341 271608
rect 114176 270843 114210 271608
rect 112367 270783 114150 270817
rect 114389 271554 115443 271588
rect 114329 270832 114363 271528
rect 115469 270832 115503 271528
rect 114389 270772 115443 270806
rect 120297 280779 121668 280813
rect 120237 269038 120271 280753
rect 121694 269038 121728 280753
rect 122238 280574 123578 280608
rect 122178 279026 122212 280548
rect 123604 279026 123638 280548
rect 122238 278966 123578 279000
rect 122314 278448 124310 278482
rect 122254 277247 122288 278422
rect 124336 277247 124370 278422
rect 122314 277187 124310 277221
rect 122374 276817 123896 276851
rect 122278 276405 122312 276755
rect 123958 276405 123992 276755
rect 122374 276309 123896 276343
rect 122379 275937 124861 275971
rect 122283 275647 122317 275875
rect 124923 275647 124957 275875
rect 122379 275551 124861 275585
rect 120297 268978 121668 269012
rect 121980 272964 123494 272998
rect 121920 269054 121954 272938
rect 123520 269054 123554 272938
rect 121980 268994 123494 269028
<< poly >>
rect 106357 280885 106489 280901
rect 106357 280851 106373 280885
rect 106473 280851 106489 280885
rect 106357 280813 106489 280851
rect 106757 280885 106889 280901
rect 106757 280851 106773 280885
rect 106873 280851 106889 280885
rect 106757 280813 106889 280851
rect 107157 280885 107289 280901
rect 107157 280851 107173 280885
rect 107273 280851 107289 280885
rect 107157 280813 107289 280851
rect 107557 280885 107689 280901
rect 107557 280851 107573 280885
rect 107673 280851 107689 280885
rect 107557 280813 107689 280851
rect 107957 280885 108089 280901
rect 107957 280851 107973 280885
rect 108073 280851 108089 280885
rect 107957 280813 108089 280851
rect 108357 280885 108489 280901
rect 108357 280851 108373 280885
rect 108473 280851 108489 280885
rect 108357 280813 108489 280851
rect 108757 280885 108889 280901
rect 108757 280851 108773 280885
rect 108873 280851 108889 280885
rect 108757 280813 108889 280851
rect 109157 280885 109289 280901
rect 109157 280851 109173 280885
rect 109273 280851 109289 280885
rect 109157 280813 109289 280851
rect 109557 280885 109689 280901
rect 109557 280851 109573 280885
rect 109673 280851 109689 280885
rect 109557 280813 109689 280851
rect 109957 280885 110089 280901
rect 109957 280851 109973 280885
rect 110073 280851 110089 280885
rect 109957 280813 110089 280851
rect 106357 279755 106489 279793
rect 106357 279721 106373 279755
rect 106473 279721 106489 279755
rect 106357 279705 106489 279721
rect 106757 279755 106889 279793
rect 106757 279721 106773 279755
rect 106873 279721 106889 279755
rect 106757 279705 106889 279721
rect 107157 279755 107289 279793
rect 107157 279721 107173 279755
rect 107273 279721 107289 279755
rect 107157 279705 107289 279721
rect 107557 279755 107689 279793
rect 107557 279721 107573 279755
rect 107673 279721 107689 279755
rect 107557 279705 107689 279721
rect 107957 279755 108089 279793
rect 107957 279721 107973 279755
rect 108073 279721 108089 279755
rect 107957 279705 108089 279721
rect 108357 279755 108489 279793
rect 108357 279721 108373 279755
rect 108473 279721 108489 279755
rect 108357 279705 108489 279721
rect 108757 279755 108889 279793
rect 108757 279721 108773 279755
rect 108873 279721 108889 279755
rect 108757 279705 108889 279721
rect 109157 279755 109289 279793
rect 109157 279721 109173 279755
rect 109273 279721 109289 279755
rect 109157 279705 109289 279721
rect 109557 279755 109689 279793
rect 109557 279721 109573 279755
rect 109673 279721 109689 279755
rect 109557 279705 109689 279721
rect 109957 279755 110089 279793
rect 109957 279721 109973 279755
rect 110073 279721 110089 279755
rect 109957 279705 110089 279721
rect 106271 278995 106368 279011
rect 106271 278773 106287 278995
rect 106321 278773 106368 278995
rect 106271 278757 106368 278773
rect 107582 278995 107679 279011
rect 107582 278773 107629 278995
rect 107663 278773 107679 278995
rect 107582 278757 107679 278773
rect 106271 278395 106368 278411
rect 106271 278173 106287 278395
rect 106321 278173 106368 278395
rect 106271 278157 106368 278173
rect 107582 278395 107679 278411
rect 107582 278173 107629 278395
rect 107663 278173 107679 278395
rect 107582 278157 107679 278173
rect 106394 277148 106491 277164
rect 106394 277106 106410 277148
rect 106444 277106 106491 277148
rect 106394 277090 106491 277106
rect 107525 277148 107622 277164
rect 107525 277106 107572 277148
rect 107606 277106 107622 277148
rect 107525 277090 107622 277106
rect 109777 279083 110063 279099
rect 109777 279049 109793 279083
rect 110047 279049 110063 279083
rect 109777 279011 110063 279049
rect 109777 277935 110063 277973
rect 109777 277901 109793 277935
rect 110047 277901 110063 277935
rect 109777 277885 110063 277901
rect 109777 277827 110063 277843
rect 109777 277793 109793 277827
rect 110047 277793 110063 277827
rect 109777 277755 110063 277793
rect 109777 276679 110063 276717
rect 109777 276645 109793 276679
rect 110047 276645 110063 276679
rect 109777 276629 110063 276645
rect 106854 275697 106951 275713
rect 106854 274951 106870 275697
rect 106904 274951 106951 275697
rect 106854 274935 106951 274951
rect 107129 275697 107226 275713
rect 107129 274951 107176 275697
rect 107210 274951 107226 275697
rect 107129 274935 107226 274951
rect 107354 275697 107451 275713
rect 107354 274951 107370 275697
rect 107404 274951 107451 275697
rect 107354 274935 107451 274951
rect 107629 275697 107726 275713
rect 107629 274951 107676 275697
rect 107710 274951 107726 275697
rect 107629 274935 107726 274951
rect 107854 275697 107951 275713
rect 107854 274951 107870 275697
rect 107904 274951 107951 275697
rect 107854 274935 107951 274951
rect 108129 275697 108226 275713
rect 108129 274951 108176 275697
rect 108210 274951 108226 275697
rect 108129 274935 108226 274951
rect 108354 275697 108451 275713
rect 108354 274951 108370 275697
rect 108404 274951 108451 275697
rect 108354 274935 108451 274951
rect 108629 275697 108726 275713
rect 108629 274951 108676 275697
rect 108710 274951 108726 275697
rect 108629 274935 108726 274951
rect 108854 275697 108951 275713
rect 108854 274951 108870 275697
rect 108904 274951 108951 275697
rect 108854 274935 108951 274951
rect 109129 275697 109226 275713
rect 109129 274951 109176 275697
rect 109210 274951 109226 275697
rect 109129 274935 109226 274951
rect 109354 275697 109451 275713
rect 109354 274951 109370 275697
rect 109404 274951 109451 275697
rect 109354 274935 109451 274951
rect 109629 275697 109726 275713
rect 109629 274951 109676 275697
rect 109710 274951 109726 275697
rect 109629 274935 109726 274951
rect 107459 272151 108079 272167
rect 107459 272117 107475 272151
rect 108063 272117 108079 272151
rect 107459 272079 108079 272117
rect 106981 272043 107191 272059
rect 106981 272009 106997 272043
rect 107175 272009 107191 272043
rect 106981 271971 107191 272009
rect 106981 271769 107191 271807
rect 106981 271735 106997 271769
rect 107175 271735 107191 271769
rect 106981 271719 107191 271735
rect 107459 271697 108079 271735
rect 107459 271663 107475 271697
rect 108063 271663 108079 271697
rect 107459 271647 108079 271663
rect 107085 271473 107173 271489
rect 107085 271327 107101 271473
rect 107135 271327 107173 271473
rect 107085 271311 107173 271327
rect 108373 271473 108461 271489
rect 108373 271327 108411 271473
rect 108445 271327 108461 271473
rect 108373 271311 108461 271327
rect 107085 271103 107173 271119
rect 107085 270957 107101 271103
rect 107135 270957 107173 271103
rect 107085 270941 107173 270957
rect 108373 271103 108461 271119
rect 108373 270957 108411 271103
rect 108445 270957 108461 271103
rect 108373 270941 108461 270957
rect 109440 272507 109510 272523
rect 109440 272473 109456 272507
rect 109494 272473 109510 272507
rect 109440 272426 109510 272473
rect 109440 270659 109510 270706
rect 109440 270625 109456 270659
rect 109494 270625 109510 270659
rect 109440 270609 109510 270625
rect 111436 280804 111524 280820
rect 111436 280676 111452 280804
rect 111486 280676 111524 280804
rect 111436 280660 111524 280676
rect 112624 280804 112712 280820
rect 112624 280676 112662 280804
rect 112696 280676 112712 280804
rect 112624 280660 112712 280676
rect 112882 280812 112970 280828
rect 112882 280644 112898 280812
rect 112932 280644 112970 280812
rect 112882 280628 112970 280644
rect 114070 280812 114158 280828
rect 114070 280644 114108 280812
rect 114142 280644 114158 280812
rect 114070 280628 114158 280644
rect 111436 280444 111524 280460
rect 111436 280316 111452 280444
rect 111486 280316 111524 280444
rect 111436 280300 111524 280316
rect 112624 280444 112712 280460
rect 112624 280316 112662 280444
rect 112696 280316 112712 280444
rect 112624 280300 112712 280316
rect 112882 280388 112970 280404
rect 112882 280220 112898 280388
rect 112932 280220 112970 280388
rect 112882 280204 112970 280220
rect 114070 280388 114158 280404
rect 114070 280220 114108 280388
rect 114142 280220 114158 280388
rect 114070 280204 114158 280220
rect 111436 280084 111524 280100
rect 111436 279956 111452 280084
rect 111486 279956 111524 280084
rect 111436 279940 111524 279956
rect 112624 280084 112712 280100
rect 112624 279956 112662 280084
rect 112696 279956 112712 280084
rect 112624 279940 112712 279956
rect 112912 279986 113000 280002
rect 112912 279938 112928 279986
rect 112962 279938 113000 279986
rect 112912 279922 113000 279938
rect 114100 279986 114188 280002
rect 114100 279938 114138 279986
rect 114172 279938 114188 279986
rect 114100 279922 114188 279938
rect 111436 279724 111524 279740
rect 111436 279596 111452 279724
rect 111486 279596 111524 279724
rect 111436 279580 111524 279596
rect 112624 279724 112712 279740
rect 112624 279596 112662 279724
rect 112696 279596 112712 279724
rect 112912 279688 113000 279704
rect 112912 279640 112928 279688
rect 112962 279640 113000 279688
rect 112912 279624 113000 279640
rect 114100 279688 114188 279704
rect 114100 279640 114138 279688
rect 114172 279640 114188 279688
rect 114100 279624 114188 279640
rect 112624 279580 112712 279596
rect 114560 280787 114657 280803
rect 114560 280419 114576 280787
rect 114610 280419 114657 280787
rect 114560 280403 114657 280419
rect 114857 280787 114954 280803
rect 114857 280419 114904 280787
rect 114938 280419 114954 280787
rect 114857 280403 114954 280419
rect 114560 280101 114657 280117
rect 114560 279973 114576 280101
rect 114610 279973 114657 280101
rect 114560 279957 114657 279973
rect 114857 280101 114954 280117
rect 114857 279973 114904 280101
rect 114938 279973 114954 280101
rect 114857 279957 114954 279973
rect 114560 279693 114657 279709
rect 114560 279565 114576 279693
rect 114610 279565 114657 279693
rect 114560 279549 114657 279565
rect 114857 279693 114954 279709
rect 114857 279565 114904 279693
rect 114938 279565 114954 279693
rect 114857 279549 114954 279565
rect 115251 280787 115348 280803
rect 115251 280419 115267 280787
rect 115301 280419 115348 280787
rect 115251 280403 115348 280419
rect 115548 280787 115645 280803
rect 115548 280419 115595 280787
rect 115629 280419 115645 280787
rect 115548 280403 115645 280419
rect 115251 280101 115348 280117
rect 115251 279973 115267 280101
rect 115301 279973 115348 280101
rect 115251 279957 115348 279973
rect 115548 280101 115645 280117
rect 115548 279973 115595 280101
rect 115629 279973 115645 280101
rect 115548 279957 115645 279973
rect 115251 279693 115348 279709
rect 115251 279565 115267 279693
rect 115301 279565 115348 279693
rect 115251 279549 115348 279565
rect 115548 279693 115645 279709
rect 115548 279565 115595 279693
rect 115629 279565 115645 279693
rect 115548 279549 115645 279565
rect 116047 280812 116135 280828
rect 116047 280644 116063 280812
rect 116097 280644 116135 280812
rect 116047 280628 116135 280644
rect 117235 280812 117323 280828
rect 117235 280644 117273 280812
rect 117307 280644 117323 280812
rect 117493 280804 117581 280820
rect 117493 280676 117509 280804
rect 117543 280676 117581 280804
rect 117493 280660 117581 280676
rect 118681 280804 118769 280820
rect 118681 280676 118719 280804
rect 118753 280676 118769 280804
rect 118681 280660 118769 280676
rect 117235 280628 117323 280644
rect 117493 280444 117581 280460
rect 116047 280388 116135 280404
rect 116047 280220 116063 280388
rect 116097 280220 116135 280388
rect 116047 280204 116135 280220
rect 117235 280388 117323 280404
rect 117235 280220 117273 280388
rect 117307 280220 117323 280388
rect 117493 280316 117509 280444
rect 117543 280316 117581 280444
rect 117493 280300 117581 280316
rect 118681 280444 118769 280460
rect 118681 280316 118719 280444
rect 118753 280316 118769 280444
rect 118681 280300 118769 280316
rect 117235 280204 117323 280220
rect 117493 280084 117581 280100
rect 116017 279986 116105 280002
rect 116017 279938 116033 279986
rect 116067 279938 116105 279986
rect 116017 279922 116105 279938
rect 117205 279986 117293 280002
rect 117205 279938 117243 279986
rect 117277 279938 117293 279986
rect 117493 279956 117509 280084
rect 117543 279956 117581 280084
rect 117493 279940 117581 279956
rect 118681 280084 118769 280100
rect 118681 279956 118719 280084
rect 118753 279956 118769 280084
rect 118681 279940 118769 279956
rect 117205 279922 117293 279938
rect 117493 279724 117581 279740
rect 116017 279688 116105 279704
rect 116017 279640 116033 279688
rect 116067 279640 116105 279688
rect 116017 279624 116105 279640
rect 117205 279688 117293 279704
rect 117205 279640 117243 279688
rect 117277 279640 117293 279688
rect 117205 279624 117293 279640
rect 117493 279596 117509 279724
rect 117543 279596 117581 279724
rect 117493 279580 117581 279596
rect 118681 279724 118769 279740
rect 118681 279596 118719 279724
rect 118753 279596 118769 279724
rect 118681 279580 118769 279596
rect 111436 279138 111524 279154
rect 111436 279010 111452 279138
rect 111486 279010 111524 279138
rect 111436 278994 111524 279010
rect 112624 279138 112712 279154
rect 112624 279010 112662 279138
rect 112696 279010 112712 279138
rect 112624 278994 112712 279010
rect 112882 279146 112970 279162
rect 112882 278978 112898 279146
rect 112932 278978 112970 279146
rect 112882 278962 112970 278978
rect 114070 279146 114158 279162
rect 114070 278978 114108 279146
rect 114142 278978 114158 279146
rect 114070 278962 114158 278978
rect 111436 278778 111524 278794
rect 111436 278650 111452 278778
rect 111486 278650 111524 278778
rect 111436 278634 111524 278650
rect 112624 278778 112712 278794
rect 112624 278650 112662 278778
rect 112696 278650 112712 278778
rect 112624 278634 112712 278650
rect 112882 278722 112970 278738
rect 112882 278554 112898 278722
rect 112932 278554 112970 278722
rect 112882 278538 112970 278554
rect 114070 278722 114158 278738
rect 114070 278554 114108 278722
rect 114142 278554 114158 278722
rect 114070 278538 114158 278554
rect 111436 278418 111524 278434
rect 111436 278290 111452 278418
rect 111486 278290 111524 278418
rect 111436 278274 111524 278290
rect 112624 278418 112712 278434
rect 112624 278290 112662 278418
rect 112696 278290 112712 278418
rect 112624 278274 112712 278290
rect 112912 278320 113000 278336
rect 112912 278272 112928 278320
rect 112962 278272 113000 278320
rect 112912 278256 113000 278272
rect 114100 278320 114188 278336
rect 114100 278272 114138 278320
rect 114172 278272 114188 278320
rect 114100 278256 114188 278272
rect 111436 278058 111524 278074
rect 111436 277930 111452 278058
rect 111486 277930 111524 278058
rect 111436 277914 111524 277930
rect 112624 278058 112712 278074
rect 112624 277930 112662 278058
rect 112696 277930 112712 278058
rect 112912 278022 113000 278038
rect 112912 277974 112928 278022
rect 112962 277974 113000 278022
rect 112912 277958 113000 277974
rect 114100 278022 114188 278038
rect 114100 277974 114138 278022
rect 114172 277974 114188 278022
rect 114100 277958 114188 277974
rect 112624 277914 112712 277930
rect 114560 279121 114657 279137
rect 114560 278753 114576 279121
rect 114610 278753 114657 279121
rect 114560 278737 114657 278753
rect 114857 279121 114954 279137
rect 114857 278753 114904 279121
rect 114938 278753 114954 279121
rect 114857 278737 114954 278753
rect 114560 278435 114657 278451
rect 114560 278307 114576 278435
rect 114610 278307 114657 278435
rect 114560 278291 114657 278307
rect 114857 278435 114954 278451
rect 114857 278307 114904 278435
rect 114938 278307 114954 278435
rect 114857 278291 114954 278307
rect 114560 278027 114657 278043
rect 114560 277899 114576 278027
rect 114610 277899 114657 278027
rect 114560 277883 114657 277899
rect 114857 278027 114954 278043
rect 114857 277899 114904 278027
rect 114938 277899 114954 278027
rect 114857 277883 114954 277899
rect 115251 279121 115348 279137
rect 115251 278753 115267 279121
rect 115301 278753 115348 279121
rect 115251 278737 115348 278753
rect 115548 279121 115645 279137
rect 115548 278753 115595 279121
rect 115629 278753 115645 279121
rect 115548 278737 115645 278753
rect 115251 278435 115348 278451
rect 115251 278307 115267 278435
rect 115301 278307 115348 278435
rect 115251 278291 115348 278307
rect 115548 278435 115645 278451
rect 115548 278307 115595 278435
rect 115629 278307 115645 278435
rect 115548 278291 115645 278307
rect 115251 278027 115348 278043
rect 115251 277899 115267 278027
rect 115301 277899 115348 278027
rect 115251 277883 115348 277899
rect 115548 278027 115645 278043
rect 115548 277899 115595 278027
rect 115629 277899 115645 278027
rect 115548 277883 115645 277899
rect 116047 279146 116135 279162
rect 116047 278978 116063 279146
rect 116097 278978 116135 279146
rect 116047 278962 116135 278978
rect 117235 279146 117323 279162
rect 117235 278978 117273 279146
rect 117307 278978 117323 279146
rect 117493 279138 117581 279154
rect 117493 279010 117509 279138
rect 117543 279010 117581 279138
rect 117493 278994 117581 279010
rect 118681 279138 118769 279154
rect 118681 279010 118719 279138
rect 118753 279010 118769 279138
rect 118681 278994 118769 279010
rect 117235 278962 117323 278978
rect 117493 278778 117581 278794
rect 116047 278722 116135 278738
rect 116047 278554 116063 278722
rect 116097 278554 116135 278722
rect 116047 278538 116135 278554
rect 117235 278722 117323 278738
rect 117235 278554 117273 278722
rect 117307 278554 117323 278722
rect 117493 278650 117509 278778
rect 117543 278650 117581 278778
rect 117493 278634 117581 278650
rect 118681 278778 118769 278794
rect 118681 278650 118719 278778
rect 118753 278650 118769 278778
rect 118681 278634 118769 278650
rect 117235 278538 117323 278554
rect 117493 278418 117581 278434
rect 116017 278320 116105 278336
rect 116017 278272 116033 278320
rect 116067 278272 116105 278320
rect 116017 278256 116105 278272
rect 117205 278320 117293 278336
rect 117205 278272 117243 278320
rect 117277 278272 117293 278320
rect 117493 278290 117509 278418
rect 117543 278290 117581 278418
rect 117493 278274 117581 278290
rect 118681 278418 118769 278434
rect 118681 278290 118719 278418
rect 118753 278290 118769 278418
rect 118681 278274 118769 278290
rect 117205 278256 117293 278272
rect 117493 278058 117581 278074
rect 116017 278022 116105 278038
rect 116017 277974 116033 278022
rect 116067 277974 116105 278022
rect 116017 277958 116105 277974
rect 117205 278022 117293 278038
rect 117205 277974 117243 278022
rect 117277 277974 117293 278022
rect 117205 277958 117293 277974
rect 117493 277930 117509 278058
rect 117543 277930 117581 278058
rect 117493 277914 117581 277930
rect 118681 278058 118769 278074
rect 118681 277930 118719 278058
rect 118753 277930 118769 278058
rect 118681 277914 118769 277930
rect 111436 277472 111524 277488
rect 111436 277344 111452 277472
rect 111486 277344 111524 277472
rect 111436 277328 111524 277344
rect 112624 277472 112712 277488
rect 112624 277344 112662 277472
rect 112696 277344 112712 277472
rect 112624 277328 112712 277344
rect 112882 277480 112970 277496
rect 112882 277312 112898 277480
rect 112932 277312 112970 277480
rect 112882 277296 112970 277312
rect 114070 277480 114158 277496
rect 114070 277312 114108 277480
rect 114142 277312 114158 277480
rect 114070 277296 114158 277312
rect 111436 277112 111524 277128
rect 111436 276984 111452 277112
rect 111486 276984 111524 277112
rect 111436 276968 111524 276984
rect 112624 277112 112712 277128
rect 112624 276984 112662 277112
rect 112696 276984 112712 277112
rect 112624 276968 112712 276984
rect 112882 277056 112970 277072
rect 112882 276888 112898 277056
rect 112932 276888 112970 277056
rect 112882 276872 112970 276888
rect 114070 277056 114158 277072
rect 114070 276888 114108 277056
rect 114142 276888 114158 277056
rect 114070 276872 114158 276888
rect 111436 276752 111524 276768
rect 111436 276624 111452 276752
rect 111486 276624 111524 276752
rect 111436 276608 111524 276624
rect 112624 276752 112712 276768
rect 112624 276624 112662 276752
rect 112696 276624 112712 276752
rect 112624 276608 112712 276624
rect 112912 276654 113000 276670
rect 112912 276606 112928 276654
rect 112962 276606 113000 276654
rect 112912 276590 113000 276606
rect 114100 276654 114188 276670
rect 114100 276606 114138 276654
rect 114172 276606 114188 276654
rect 114100 276590 114188 276606
rect 111436 276392 111524 276408
rect 111436 276264 111452 276392
rect 111486 276264 111524 276392
rect 111436 276248 111524 276264
rect 112624 276392 112712 276408
rect 112624 276264 112662 276392
rect 112696 276264 112712 276392
rect 112912 276356 113000 276372
rect 112912 276308 112928 276356
rect 112962 276308 113000 276356
rect 112912 276292 113000 276308
rect 114100 276356 114188 276372
rect 114100 276308 114138 276356
rect 114172 276308 114188 276356
rect 114100 276292 114188 276308
rect 112624 276248 112712 276264
rect 114560 277455 114657 277471
rect 114560 277087 114576 277455
rect 114610 277087 114657 277455
rect 114560 277071 114657 277087
rect 114857 277455 114954 277471
rect 114857 277087 114904 277455
rect 114938 277087 114954 277455
rect 114857 277071 114954 277087
rect 114560 276769 114657 276785
rect 114560 276641 114576 276769
rect 114610 276641 114657 276769
rect 114560 276625 114657 276641
rect 114857 276769 114954 276785
rect 114857 276641 114904 276769
rect 114938 276641 114954 276769
rect 114857 276625 114954 276641
rect 114560 276361 114657 276377
rect 114560 276233 114576 276361
rect 114610 276233 114657 276361
rect 114560 276217 114657 276233
rect 114857 276361 114954 276377
rect 114857 276233 114904 276361
rect 114938 276233 114954 276361
rect 114857 276217 114954 276233
rect 115251 277455 115348 277471
rect 115251 277087 115267 277455
rect 115301 277087 115348 277455
rect 115251 277071 115348 277087
rect 115548 277455 115645 277471
rect 115548 277087 115595 277455
rect 115629 277087 115645 277455
rect 115548 277071 115645 277087
rect 115251 276769 115348 276785
rect 115251 276641 115267 276769
rect 115301 276641 115348 276769
rect 115251 276625 115348 276641
rect 115548 276769 115645 276785
rect 115548 276641 115595 276769
rect 115629 276641 115645 276769
rect 115548 276625 115645 276641
rect 115251 276361 115348 276377
rect 115251 276233 115267 276361
rect 115301 276233 115348 276361
rect 115251 276217 115348 276233
rect 115548 276361 115645 276377
rect 115548 276233 115595 276361
rect 115629 276233 115645 276361
rect 115548 276217 115645 276233
rect 116047 277480 116135 277496
rect 116047 277312 116063 277480
rect 116097 277312 116135 277480
rect 116047 277296 116135 277312
rect 117235 277480 117323 277496
rect 117235 277312 117273 277480
rect 117307 277312 117323 277480
rect 117493 277472 117581 277488
rect 117493 277344 117509 277472
rect 117543 277344 117581 277472
rect 117493 277328 117581 277344
rect 118681 277472 118769 277488
rect 118681 277344 118719 277472
rect 118753 277344 118769 277472
rect 118681 277328 118769 277344
rect 117235 277296 117323 277312
rect 117493 277112 117581 277128
rect 116047 277056 116135 277072
rect 116047 276888 116063 277056
rect 116097 276888 116135 277056
rect 116047 276872 116135 276888
rect 117235 277056 117323 277072
rect 117235 276888 117273 277056
rect 117307 276888 117323 277056
rect 117493 276984 117509 277112
rect 117543 276984 117581 277112
rect 117493 276968 117581 276984
rect 118681 277112 118769 277128
rect 118681 276984 118719 277112
rect 118753 276984 118769 277112
rect 118681 276968 118769 276984
rect 117235 276872 117323 276888
rect 117493 276752 117581 276768
rect 116017 276654 116105 276670
rect 116017 276606 116033 276654
rect 116067 276606 116105 276654
rect 116017 276590 116105 276606
rect 117205 276654 117293 276670
rect 117205 276606 117243 276654
rect 117277 276606 117293 276654
rect 117493 276624 117509 276752
rect 117543 276624 117581 276752
rect 117493 276608 117581 276624
rect 118681 276752 118769 276768
rect 118681 276624 118719 276752
rect 118753 276624 118769 276752
rect 118681 276608 118769 276624
rect 117205 276590 117293 276606
rect 117493 276392 117581 276408
rect 116017 276356 116105 276372
rect 116017 276308 116033 276356
rect 116067 276308 116105 276356
rect 116017 276292 116105 276308
rect 117205 276356 117293 276372
rect 117205 276308 117243 276356
rect 117277 276308 117293 276356
rect 117205 276292 117293 276308
rect 117493 276264 117509 276392
rect 117543 276264 117581 276392
rect 117493 276248 117581 276264
rect 118681 276392 118769 276408
rect 118681 276264 118719 276392
rect 118753 276264 118769 276392
rect 118681 276248 118769 276264
rect 111436 275806 111524 275822
rect 111436 275678 111452 275806
rect 111486 275678 111524 275806
rect 111436 275662 111524 275678
rect 112624 275806 112712 275822
rect 112624 275678 112662 275806
rect 112696 275678 112712 275806
rect 112624 275662 112712 275678
rect 112882 275814 112970 275830
rect 112882 275646 112898 275814
rect 112932 275646 112970 275814
rect 112882 275630 112970 275646
rect 114070 275814 114158 275830
rect 114070 275646 114108 275814
rect 114142 275646 114158 275814
rect 114070 275630 114158 275646
rect 111436 275446 111524 275462
rect 111436 275318 111452 275446
rect 111486 275318 111524 275446
rect 111436 275302 111524 275318
rect 112624 275446 112712 275462
rect 112624 275318 112662 275446
rect 112696 275318 112712 275446
rect 112624 275302 112712 275318
rect 112882 275390 112970 275406
rect 112882 275222 112898 275390
rect 112932 275222 112970 275390
rect 112882 275206 112970 275222
rect 114070 275390 114158 275406
rect 114070 275222 114108 275390
rect 114142 275222 114158 275390
rect 114070 275206 114158 275222
rect 111436 275086 111524 275102
rect 111436 274958 111452 275086
rect 111486 274958 111524 275086
rect 111436 274942 111524 274958
rect 112624 275086 112712 275102
rect 112624 274958 112662 275086
rect 112696 274958 112712 275086
rect 112624 274942 112712 274958
rect 112912 274988 113000 275004
rect 112912 274940 112928 274988
rect 112962 274940 113000 274988
rect 112912 274924 113000 274940
rect 114100 274988 114188 275004
rect 114100 274940 114138 274988
rect 114172 274940 114188 274988
rect 114100 274924 114188 274940
rect 111436 274726 111524 274742
rect 111436 274598 111452 274726
rect 111486 274598 111524 274726
rect 111436 274582 111524 274598
rect 112624 274726 112712 274742
rect 112624 274598 112662 274726
rect 112696 274598 112712 274726
rect 112912 274690 113000 274706
rect 112912 274642 112928 274690
rect 112962 274642 113000 274690
rect 112912 274626 113000 274642
rect 114100 274690 114188 274706
rect 114100 274642 114138 274690
rect 114172 274642 114188 274690
rect 114100 274626 114188 274642
rect 112624 274582 112712 274598
rect 114560 275789 114657 275805
rect 114560 275421 114576 275789
rect 114610 275421 114657 275789
rect 114560 275405 114657 275421
rect 114857 275789 114954 275805
rect 114857 275421 114904 275789
rect 114938 275421 114954 275789
rect 114857 275405 114954 275421
rect 114560 275103 114657 275119
rect 114560 274975 114576 275103
rect 114610 274975 114657 275103
rect 114560 274959 114657 274975
rect 114857 275103 114954 275119
rect 114857 274975 114904 275103
rect 114938 274975 114954 275103
rect 114857 274959 114954 274975
rect 114560 274695 114657 274711
rect 114560 274567 114576 274695
rect 114610 274567 114657 274695
rect 114560 274551 114657 274567
rect 114857 274695 114954 274711
rect 114857 274567 114904 274695
rect 114938 274567 114954 274695
rect 114857 274551 114954 274567
rect 115251 275789 115348 275805
rect 115251 275421 115267 275789
rect 115301 275421 115348 275789
rect 115251 275405 115348 275421
rect 115548 275789 115645 275805
rect 115548 275421 115595 275789
rect 115629 275421 115645 275789
rect 115548 275405 115645 275421
rect 115251 275103 115348 275119
rect 115251 274975 115267 275103
rect 115301 274975 115348 275103
rect 115251 274959 115348 274975
rect 115548 275103 115645 275119
rect 115548 274975 115595 275103
rect 115629 274975 115645 275103
rect 115548 274959 115645 274975
rect 115251 274695 115348 274711
rect 115251 274567 115267 274695
rect 115301 274567 115348 274695
rect 115251 274551 115348 274567
rect 115548 274695 115645 274711
rect 115548 274567 115595 274695
rect 115629 274567 115645 274695
rect 115548 274551 115645 274567
rect 116047 275814 116135 275830
rect 116047 275646 116063 275814
rect 116097 275646 116135 275814
rect 116047 275630 116135 275646
rect 117235 275814 117323 275830
rect 117235 275646 117273 275814
rect 117307 275646 117323 275814
rect 117493 275806 117581 275822
rect 117493 275678 117509 275806
rect 117543 275678 117581 275806
rect 117493 275662 117581 275678
rect 118681 275806 118769 275822
rect 118681 275678 118719 275806
rect 118753 275678 118769 275806
rect 118681 275662 118769 275678
rect 117235 275630 117323 275646
rect 117493 275446 117581 275462
rect 116047 275390 116135 275406
rect 116047 275222 116063 275390
rect 116097 275222 116135 275390
rect 116047 275206 116135 275222
rect 117235 275390 117323 275406
rect 117235 275222 117273 275390
rect 117307 275222 117323 275390
rect 117493 275318 117509 275446
rect 117543 275318 117581 275446
rect 117493 275302 117581 275318
rect 118681 275446 118769 275462
rect 118681 275318 118719 275446
rect 118753 275318 118769 275446
rect 118681 275302 118769 275318
rect 117235 275206 117323 275222
rect 117493 275086 117581 275102
rect 116017 274988 116105 275004
rect 116017 274940 116033 274988
rect 116067 274940 116105 274988
rect 116017 274924 116105 274940
rect 117205 274988 117293 275004
rect 117205 274940 117243 274988
rect 117277 274940 117293 274988
rect 117493 274958 117509 275086
rect 117543 274958 117581 275086
rect 117493 274942 117581 274958
rect 118681 275086 118769 275102
rect 118681 274958 118719 275086
rect 118753 274958 118769 275086
rect 118681 274942 118769 274958
rect 117205 274924 117293 274940
rect 117493 274726 117581 274742
rect 116017 274690 116105 274706
rect 116017 274642 116033 274690
rect 116067 274642 116105 274690
rect 116017 274626 116105 274642
rect 117205 274690 117293 274706
rect 117205 274642 117243 274690
rect 117277 274642 117293 274690
rect 117205 274626 117293 274642
rect 117493 274598 117509 274726
rect 117543 274598 117581 274726
rect 117493 274582 117581 274598
rect 118681 274726 118769 274742
rect 118681 274598 118719 274726
rect 118753 274598 118769 274726
rect 118681 274582 118769 274598
rect 111436 274140 111524 274156
rect 111436 274012 111452 274140
rect 111486 274012 111524 274140
rect 111436 273996 111524 274012
rect 112624 274140 112712 274156
rect 112624 274012 112662 274140
rect 112696 274012 112712 274140
rect 112624 273996 112712 274012
rect 112882 274148 112970 274164
rect 112882 273980 112898 274148
rect 112932 273980 112970 274148
rect 112882 273964 112970 273980
rect 114070 274148 114158 274164
rect 114070 273980 114108 274148
rect 114142 273980 114158 274148
rect 114070 273964 114158 273980
rect 111436 273780 111524 273796
rect 111436 273652 111452 273780
rect 111486 273652 111524 273780
rect 111436 273636 111524 273652
rect 112624 273780 112712 273796
rect 112624 273652 112662 273780
rect 112696 273652 112712 273780
rect 112624 273636 112712 273652
rect 112882 273724 112970 273740
rect 112882 273556 112898 273724
rect 112932 273556 112970 273724
rect 112882 273540 112970 273556
rect 114070 273724 114158 273740
rect 114070 273556 114108 273724
rect 114142 273556 114158 273724
rect 114070 273540 114158 273556
rect 111436 273420 111524 273436
rect 111436 273292 111452 273420
rect 111486 273292 111524 273420
rect 111436 273276 111524 273292
rect 112624 273420 112712 273436
rect 112624 273292 112662 273420
rect 112696 273292 112712 273420
rect 112624 273276 112712 273292
rect 112912 273322 113000 273338
rect 112912 273274 112928 273322
rect 112962 273274 113000 273322
rect 112912 273258 113000 273274
rect 114100 273322 114188 273338
rect 114100 273274 114138 273322
rect 114172 273274 114188 273322
rect 114100 273258 114188 273274
rect 111436 273060 111524 273076
rect 111436 272932 111452 273060
rect 111486 272932 111524 273060
rect 111436 272916 111524 272932
rect 112624 273060 112712 273076
rect 112624 272932 112662 273060
rect 112696 272932 112712 273060
rect 112912 273024 113000 273040
rect 112912 272976 112928 273024
rect 112962 272976 113000 273024
rect 112912 272960 113000 272976
rect 114100 273024 114188 273040
rect 114100 272976 114138 273024
rect 114172 272976 114188 273024
rect 114100 272960 114188 272976
rect 112624 272916 112712 272932
rect 114560 274123 114657 274139
rect 114560 273755 114576 274123
rect 114610 273755 114657 274123
rect 114560 273739 114657 273755
rect 114857 274123 114954 274139
rect 114857 273755 114904 274123
rect 114938 273755 114954 274123
rect 114857 273739 114954 273755
rect 114560 273437 114657 273453
rect 114560 273309 114576 273437
rect 114610 273309 114657 273437
rect 114560 273293 114657 273309
rect 114857 273437 114954 273453
rect 114857 273309 114904 273437
rect 114938 273309 114954 273437
rect 114857 273293 114954 273309
rect 114560 273029 114657 273045
rect 114560 272901 114576 273029
rect 114610 272901 114657 273029
rect 114560 272885 114657 272901
rect 114857 273029 114954 273045
rect 114857 272901 114904 273029
rect 114938 272901 114954 273029
rect 114857 272885 114954 272901
rect 115251 274123 115348 274139
rect 115251 273755 115267 274123
rect 115301 273755 115348 274123
rect 115251 273739 115348 273755
rect 115548 274123 115645 274139
rect 115548 273755 115595 274123
rect 115629 273755 115645 274123
rect 115548 273739 115645 273755
rect 115251 273437 115348 273453
rect 115251 273309 115267 273437
rect 115301 273309 115348 273437
rect 115251 273293 115348 273309
rect 115548 273437 115645 273453
rect 115548 273309 115595 273437
rect 115629 273309 115645 273437
rect 115548 273293 115645 273309
rect 115251 273029 115348 273045
rect 115251 272901 115267 273029
rect 115301 272901 115348 273029
rect 115251 272885 115348 272901
rect 115548 273029 115645 273045
rect 115548 272901 115595 273029
rect 115629 272901 115645 273029
rect 115548 272885 115645 272901
rect 116047 274148 116135 274164
rect 116047 273980 116063 274148
rect 116097 273980 116135 274148
rect 116047 273964 116135 273980
rect 117235 274148 117323 274164
rect 117235 273980 117273 274148
rect 117307 273980 117323 274148
rect 117493 274140 117581 274156
rect 117493 274012 117509 274140
rect 117543 274012 117581 274140
rect 117493 273996 117581 274012
rect 118681 274140 118769 274156
rect 118681 274012 118719 274140
rect 118753 274012 118769 274140
rect 118681 273996 118769 274012
rect 117235 273964 117323 273980
rect 117493 273780 117581 273796
rect 116047 273724 116135 273740
rect 116047 273556 116063 273724
rect 116097 273556 116135 273724
rect 116047 273540 116135 273556
rect 117235 273724 117323 273740
rect 117235 273556 117273 273724
rect 117307 273556 117323 273724
rect 117493 273652 117509 273780
rect 117543 273652 117581 273780
rect 117493 273636 117581 273652
rect 118681 273780 118769 273796
rect 118681 273652 118719 273780
rect 118753 273652 118769 273780
rect 118681 273636 118769 273652
rect 117235 273540 117323 273556
rect 117493 273420 117581 273436
rect 116017 273322 116105 273338
rect 116017 273274 116033 273322
rect 116067 273274 116105 273322
rect 116017 273258 116105 273274
rect 117205 273322 117293 273338
rect 117205 273274 117243 273322
rect 117277 273274 117293 273322
rect 117493 273292 117509 273420
rect 117543 273292 117581 273420
rect 117493 273276 117581 273292
rect 118681 273420 118769 273436
rect 118681 273292 118719 273420
rect 118753 273292 118769 273420
rect 118681 273276 118769 273292
rect 117205 273258 117293 273274
rect 117493 273060 117581 273076
rect 116017 273024 116105 273040
rect 116017 272976 116033 273024
rect 116067 272976 116105 273024
rect 116017 272960 116105 272976
rect 117205 273024 117293 273040
rect 117205 272976 117243 273024
rect 117277 272976 117293 273024
rect 117205 272960 117293 272976
rect 117493 272932 117509 273060
rect 117543 272932 117581 273060
rect 117493 272916 117581 272932
rect 118681 273060 118769 273076
rect 118681 272932 118719 273060
rect 118753 272932 118769 273060
rect 118681 272916 118769 272932
rect 115881 271996 116041 272012
rect 115881 271962 115897 271996
rect 116025 271962 116041 271996
rect 115881 271924 116041 271962
rect 116281 271996 116441 272012
rect 116281 271962 116297 271996
rect 116425 271962 116441 271996
rect 116281 271924 116441 271962
rect 116681 271996 116841 272012
rect 116681 271962 116697 271996
rect 116825 271962 116841 271996
rect 116681 271924 116841 271962
rect 117081 271996 117241 272012
rect 117081 271962 117097 271996
rect 117225 271962 117241 271996
rect 117081 271924 117241 271962
rect 117481 271996 117641 272012
rect 117481 271962 117497 271996
rect 117625 271962 117641 271996
rect 117481 271924 117641 271962
rect 117881 271996 118041 272012
rect 117881 271962 117897 271996
rect 118025 271962 118041 271996
rect 117881 271924 118041 271962
rect 118281 271996 118441 272012
rect 118281 271962 118297 271996
rect 118425 271962 118441 271996
rect 118281 271924 118441 271962
rect 118681 271996 118841 272012
rect 118681 271962 118697 271996
rect 118825 271962 118841 271996
rect 118681 271924 118841 271962
rect 112578 271387 112738 271403
rect 112578 271353 112594 271387
rect 112722 271353 112738 271387
rect 112578 271306 112738 271353
rect 112978 271387 113138 271403
rect 112978 271353 112994 271387
rect 113122 271353 113138 271387
rect 112978 271306 113138 271353
rect 113378 271387 113538 271403
rect 113378 271353 113394 271387
rect 113522 271353 113538 271387
rect 113378 271306 113538 271353
rect 113778 271387 113938 271403
rect 113778 271353 113794 271387
rect 113922 271353 113938 271387
rect 113778 271306 113938 271353
rect 112578 271059 112738 271106
rect 112578 271025 112594 271059
rect 112722 271025 112738 271059
rect 112578 271009 112738 271025
rect 112978 271059 113138 271106
rect 112978 271025 112994 271059
rect 113122 271025 113138 271059
rect 112978 271009 113138 271025
rect 113378 271059 113538 271106
rect 113378 271025 113394 271059
rect 113522 271025 113538 271059
rect 113378 271009 113538 271025
rect 113778 271059 113938 271106
rect 113778 271025 113794 271059
rect 113922 271025 113938 271059
rect 113778 271009 113938 271025
rect 114637 271358 114797 271374
rect 114637 271324 114653 271358
rect 114781 271324 114797 271358
rect 114637 271277 114797 271324
rect 115037 271358 115197 271374
rect 115037 271324 115053 271358
rect 115181 271324 115197 271358
rect 115037 271277 115197 271324
rect 114637 271030 114797 271077
rect 114637 270996 114653 271030
rect 114781 270996 114797 271030
rect 114637 270980 114797 270996
rect 115037 271030 115197 271077
rect 115037 270996 115053 271030
rect 115181 270996 115197 271030
rect 115037 270980 115197 270996
rect 115881 270786 116041 270824
rect 115881 270752 115897 270786
rect 116025 270752 116041 270786
rect 115881 270736 116041 270752
rect 116281 270786 116441 270824
rect 116281 270752 116297 270786
rect 116425 270752 116441 270786
rect 116281 270736 116441 270752
rect 116681 270786 116841 270824
rect 116681 270752 116697 270786
rect 116825 270752 116841 270786
rect 116681 270736 116841 270752
rect 117081 270786 117241 270824
rect 117081 270752 117097 270786
rect 117225 270752 117241 270786
rect 117081 270736 117241 270752
rect 117481 270786 117641 270824
rect 117481 270752 117497 270786
rect 117625 270752 117641 270786
rect 117481 270736 117641 270752
rect 117881 270786 118041 270824
rect 117881 270752 117897 270786
rect 118025 270752 118041 270786
rect 117881 270736 118041 270752
rect 118281 270786 118441 270824
rect 118281 270752 118297 270786
rect 118425 270752 118441 270786
rect 118281 270736 118441 270752
rect 118681 270786 118841 270824
rect 118681 270752 118697 270786
rect 118825 270752 118841 270786
rect 118681 270736 118841 270752
rect 112560 270296 112720 270312
rect 112560 270262 112576 270296
rect 112704 270262 112720 270296
rect 112560 270224 112720 270262
rect 112960 270296 113120 270312
rect 112960 270262 112976 270296
rect 113104 270262 113120 270296
rect 112960 270224 113120 270262
rect 113360 270296 113520 270312
rect 113360 270262 113376 270296
rect 113504 270262 113520 270296
rect 113360 270224 113520 270262
rect 113760 270296 113920 270312
rect 113760 270262 113776 270296
rect 113904 270262 113920 270296
rect 113760 270224 113920 270262
rect 114160 270296 114320 270312
rect 114160 270262 114176 270296
rect 114304 270262 114320 270296
rect 114160 270224 114320 270262
rect 114560 270296 114720 270312
rect 114560 270262 114576 270296
rect 114704 270262 114720 270296
rect 114560 270224 114720 270262
rect 114960 270296 115120 270312
rect 114960 270262 114976 270296
rect 115104 270262 115120 270296
rect 114960 270224 115120 270262
rect 115360 270296 115520 270312
rect 115360 270262 115376 270296
rect 115504 270262 115520 270296
rect 115360 270224 115520 270262
rect 115760 270296 115920 270312
rect 115760 270262 115776 270296
rect 115904 270262 115920 270296
rect 115760 270224 115920 270262
rect 116160 270296 116320 270312
rect 116160 270262 116176 270296
rect 116304 270262 116320 270296
rect 116160 270224 116320 270262
rect 116560 270296 116720 270312
rect 116560 270262 116576 270296
rect 116704 270262 116720 270296
rect 116560 270224 116720 270262
rect 116960 270296 117120 270312
rect 116960 270262 116976 270296
rect 117104 270262 117120 270296
rect 116960 270224 117120 270262
rect 117360 270296 117520 270312
rect 117360 270262 117376 270296
rect 117504 270262 117520 270296
rect 117360 270224 117520 270262
rect 117760 270296 117920 270312
rect 117760 270262 117776 270296
rect 117904 270262 117920 270296
rect 117760 270224 117920 270262
rect 118160 270296 118320 270312
rect 118160 270262 118176 270296
rect 118304 270262 118320 270296
rect 118160 270224 118320 270262
rect 118560 270296 118720 270312
rect 118560 270262 118576 270296
rect 118704 270262 118720 270296
rect 118560 270224 118720 270262
rect 112560 269086 112720 269124
rect 112560 269052 112576 269086
rect 112704 269052 112720 269086
rect 112560 269036 112720 269052
rect 112960 269086 113120 269124
rect 112960 269052 112976 269086
rect 113104 269052 113120 269086
rect 112960 269036 113120 269052
rect 113360 269086 113520 269124
rect 113360 269052 113376 269086
rect 113504 269052 113520 269086
rect 113360 269036 113520 269052
rect 113760 269086 113920 269124
rect 113760 269052 113776 269086
rect 113904 269052 113920 269086
rect 113760 269036 113920 269052
rect 114160 269086 114320 269124
rect 114160 269052 114176 269086
rect 114304 269052 114320 269086
rect 114160 269036 114320 269052
rect 114560 269086 114720 269124
rect 114560 269052 114576 269086
rect 114704 269052 114720 269086
rect 114560 269036 114720 269052
rect 114960 269086 115120 269124
rect 114960 269052 114976 269086
rect 115104 269052 115120 269086
rect 114960 269036 115120 269052
rect 115360 269086 115520 269124
rect 115360 269052 115376 269086
rect 115504 269052 115520 269086
rect 115360 269036 115520 269052
rect 115760 269086 115920 269124
rect 115760 269052 115776 269086
rect 115904 269052 115920 269086
rect 115760 269036 115920 269052
rect 116160 269086 116320 269124
rect 116160 269052 116176 269086
rect 116304 269052 116320 269086
rect 116160 269036 116320 269052
rect 116560 269086 116720 269124
rect 116560 269052 116576 269086
rect 116704 269052 116720 269086
rect 116560 269036 116720 269052
rect 116960 269086 117120 269124
rect 116960 269052 116976 269086
rect 117104 269052 117120 269086
rect 116960 269036 117120 269052
rect 117360 269086 117520 269124
rect 117360 269052 117376 269086
rect 117504 269052 117520 269086
rect 117360 269036 117520 269052
rect 117760 269086 117920 269124
rect 117760 269052 117776 269086
rect 117904 269052 117920 269086
rect 117760 269036 117920 269052
rect 118160 269086 118320 269124
rect 118160 269052 118176 269086
rect 118304 269052 118320 269086
rect 118160 269036 118320 269052
rect 118560 269086 118720 269124
rect 118560 269052 118576 269086
rect 118704 269052 118720 269086
rect 118560 269036 118720 269052
rect 120429 280718 120829 280734
rect 120429 280684 120445 280718
rect 120813 280684 120829 280718
rect 120429 280637 120829 280684
rect 121129 280718 121529 280734
rect 121129 280684 121145 280718
rect 121513 280684 121529 280718
rect 121129 280637 121529 280684
rect 120429 280490 120829 280537
rect 120429 280456 120445 280490
rect 120813 280456 120829 280490
rect 120429 280440 120829 280456
rect 121129 280490 121529 280537
rect 121129 280456 121145 280490
rect 121513 280456 121529 280490
rect 121129 280440 121529 280456
rect 120429 280334 120829 280350
rect 120429 280300 120445 280334
rect 120813 280300 120829 280334
rect 120429 280253 120829 280300
rect 121129 280334 121529 280350
rect 121129 280300 121145 280334
rect 121513 280300 121529 280334
rect 121129 280253 121529 280300
rect 120429 279706 120829 279753
rect 120429 279672 120445 279706
rect 120813 279672 120829 279706
rect 120429 279656 120829 279672
rect 121129 279706 121529 279753
rect 121129 279672 121145 279706
rect 121513 279672 121529 279706
rect 121129 279656 121529 279672
rect 120429 279550 120829 279566
rect 120429 279516 120445 279550
rect 120813 279516 120829 279550
rect 120429 279469 120829 279516
rect 121129 279550 121529 279566
rect 121129 279516 121145 279550
rect 121513 279516 121529 279550
rect 121129 279469 121529 279516
rect 120429 278922 120829 278969
rect 120429 278888 120445 278922
rect 120813 278888 120829 278922
rect 120429 278872 120829 278888
rect 121129 278922 121529 278969
rect 121129 278888 121145 278922
rect 121513 278888 121529 278922
rect 121129 278872 121529 278888
rect 120429 278766 120829 278782
rect 120429 278732 120445 278766
rect 120813 278732 120829 278766
rect 120429 278685 120829 278732
rect 121129 278766 121529 278782
rect 121129 278732 121145 278766
rect 121513 278732 121529 278766
rect 121129 278685 121529 278732
rect 120429 278138 120829 278185
rect 120429 278104 120445 278138
rect 120813 278104 120829 278138
rect 120429 278088 120829 278104
rect 121129 278138 121529 278185
rect 121129 278104 121145 278138
rect 121513 278104 121529 278138
rect 121129 278088 121529 278104
rect 120429 277982 120829 277998
rect 120429 277948 120445 277982
rect 120813 277948 120829 277982
rect 120429 277901 120829 277948
rect 121129 277982 121529 277998
rect 121129 277948 121145 277982
rect 121513 277948 121529 277982
rect 121129 277901 121529 277948
rect 120429 277354 120829 277401
rect 120429 277320 120445 277354
rect 120813 277320 120829 277354
rect 120429 277304 120829 277320
rect 121129 277354 121529 277401
rect 121129 277320 121145 277354
rect 121513 277320 121529 277354
rect 121129 277304 121529 277320
rect 120429 277198 120829 277214
rect 120429 277164 120445 277198
rect 120813 277164 120829 277198
rect 120429 277117 120829 277164
rect 121129 277198 121529 277214
rect 121129 277164 121145 277198
rect 121513 277164 121529 277198
rect 121129 277117 121529 277164
rect 120429 276570 120829 276617
rect 120429 276536 120445 276570
rect 120813 276536 120829 276570
rect 120429 276520 120829 276536
rect 121129 276570 121529 276617
rect 121129 276536 121145 276570
rect 121513 276536 121529 276570
rect 121129 276520 121529 276536
rect 120429 276414 120829 276430
rect 120429 276380 120445 276414
rect 120813 276380 120829 276414
rect 120429 276333 120829 276380
rect 121129 276414 121529 276430
rect 121129 276380 121145 276414
rect 121513 276380 121529 276414
rect 121129 276333 121529 276380
rect 120429 275786 120829 275833
rect 120429 275752 120445 275786
rect 120813 275752 120829 275786
rect 120429 275736 120829 275752
rect 121129 275786 121529 275833
rect 121129 275752 121145 275786
rect 121513 275752 121529 275786
rect 121129 275736 121529 275752
rect 120429 275630 120829 275646
rect 120429 275596 120445 275630
rect 120813 275596 120829 275630
rect 120429 275549 120829 275596
rect 121129 275630 121529 275646
rect 121129 275596 121145 275630
rect 121513 275596 121529 275630
rect 121129 275549 121529 275596
rect 120429 275002 120829 275049
rect 120429 274968 120445 275002
rect 120813 274968 120829 275002
rect 120429 274952 120829 274968
rect 121129 275002 121529 275049
rect 121129 274968 121145 275002
rect 121513 274968 121529 275002
rect 121129 274952 121529 274968
rect 120429 274846 120829 274862
rect 120429 274812 120445 274846
rect 120813 274812 120829 274846
rect 120429 274765 120829 274812
rect 121129 274846 121529 274862
rect 121129 274812 121145 274846
rect 121513 274812 121529 274846
rect 121129 274765 121529 274812
rect 120429 274218 120829 274265
rect 120429 274184 120445 274218
rect 120813 274184 120829 274218
rect 120429 274168 120829 274184
rect 121129 274218 121529 274265
rect 121129 274184 121145 274218
rect 121513 274184 121529 274218
rect 121129 274168 121529 274184
rect 120429 274062 120829 274078
rect 120429 274028 120445 274062
rect 120813 274028 120829 274062
rect 120429 273981 120829 274028
rect 121129 274062 121529 274078
rect 121129 274028 121145 274062
rect 121513 274028 121529 274062
rect 121129 273981 121529 274028
rect 120429 273434 120829 273481
rect 120429 273400 120445 273434
rect 120813 273400 120829 273434
rect 120429 273384 120829 273400
rect 121129 273434 121529 273481
rect 121129 273400 121145 273434
rect 121513 273400 121529 273434
rect 121129 273384 121529 273400
rect 120429 273278 120829 273294
rect 120429 273244 120445 273278
rect 120813 273244 120829 273278
rect 120429 273197 120829 273244
rect 121129 273278 121529 273294
rect 121129 273244 121145 273278
rect 121513 273244 121529 273278
rect 121129 273197 121529 273244
rect 120429 272650 120829 272697
rect 120429 272616 120445 272650
rect 120813 272616 120829 272650
rect 120429 272600 120829 272616
rect 121129 272650 121529 272697
rect 121129 272616 121145 272650
rect 121513 272616 121529 272650
rect 121129 272600 121529 272616
rect 120429 272494 120829 272510
rect 120429 272460 120445 272494
rect 120813 272460 120829 272494
rect 120429 272413 120829 272460
rect 121129 272494 121529 272510
rect 121129 272460 121145 272494
rect 121513 272460 121529 272494
rect 121129 272413 121529 272460
rect 120429 271866 120829 271913
rect 120429 271832 120445 271866
rect 120813 271832 120829 271866
rect 120429 271816 120829 271832
rect 121129 271866 121529 271913
rect 121129 271832 121145 271866
rect 121513 271832 121529 271866
rect 121129 271816 121529 271832
rect 120429 271710 120829 271726
rect 120429 271676 120445 271710
rect 120813 271676 120829 271710
rect 120429 271629 120829 271676
rect 121129 271710 121529 271726
rect 121129 271676 121145 271710
rect 121513 271676 121529 271710
rect 121129 271629 121529 271676
rect 120429 271082 120829 271129
rect 120429 271048 120445 271082
rect 120813 271048 120829 271082
rect 120429 271032 120829 271048
rect 121129 271082 121529 271129
rect 121129 271048 121145 271082
rect 121513 271048 121529 271082
rect 121129 271032 121529 271048
rect 120429 270926 120829 270942
rect 120429 270892 120445 270926
rect 120813 270892 120829 270926
rect 120429 270845 120829 270892
rect 121129 270926 121529 270942
rect 121129 270892 121145 270926
rect 121513 270892 121529 270926
rect 121129 270845 121529 270892
rect 120429 270298 120829 270345
rect 120429 270264 120445 270298
rect 120813 270264 120829 270298
rect 120429 270248 120829 270264
rect 121129 270298 121529 270345
rect 121129 270264 121145 270298
rect 121513 270264 121529 270298
rect 121129 270248 121529 270264
rect 120429 270142 120829 270158
rect 120429 270108 120445 270142
rect 120813 270108 120829 270142
rect 120429 270061 120829 270108
rect 121129 270142 121529 270158
rect 121129 270108 121145 270142
rect 121513 270108 121529 270142
rect 121129 270061 121529 270108
rect 120429 269514 120829 269561
rect 120429 269480 120445 269514
rect 120813 269480 120829 269514
rect 120429 269464 120829 269480
rect 121129 269514 121529 269561
rect 121129 269480 121145 269514
rect 121513 269480 121529 269514
rect 121129 269464 121529 269480
rect 120429 269358 120829 269374
rect 120429 269324 120445 269358
rect 120813 269324 120829 269358
rect 120429 269277 120829 269324
rect 121129 269358 121529 269374
rect 121129 269324 121145 269358
rect 121513 269324 121529 269358
rect 121129 269277 121529 269324
rect 120429 269130 120829 269177
rect 120429 269096 120445 269130
rect 120813 269096 120829 269130
rect 120429 269080 120829 269096
rect 121129 269130 121529 269177
rect 121129 269096 121145 269130
rect 121513 269096 121529 269130
rect 121129 269080 121529 269096
rect 122356 280504 122756 280520
rect 122356 280470 122372 280504
rect 122740 280470 122756 280504
rect 122356 280423 122756 280470
rect 123056 280504 123456 280520
rect 123056 280470 123072 280504
rect 123440 280470 123456 280504
rect 123056 280423 123456 280470
rect 122356 279876 122756 279923
rect 122356 279842 122372 279876
rect 122740 279842 122756 279876
rect 122356 279826 122756 279842
rect 123056 279876 123456 279923
rect 123056 279842 123072 279876
rect 123440 279842 123456 279876
rect 123056 279826 123456 279842
rect 122356 279720 122756 279736
rect 122356 279686 122372 279720
rect 122740 279686 122756 279720
rect 122356 279639 122756 279686
rect 123056 279720 123456 279736
rect 123056 279686 123072 279720
rect 123440 279686 123456 279720
rect 123056 279639 123456 279686
rect 122356 279092 122756 279139
rect 122356 279058 122372 279092
rect 122740 279058 122756 279092
rect 122356 279042 122756 279058
rect 123056 279092 123456 279139
rect 123056 279058 123072 279092
rect 123440 279058 123456 279092
rect 123056 279042 123456 279058
rect 122414 278347 123290 278363
rect 122414 278313 122430 278347
rect 123274 278313 123290 278347
rect 122414 278266 123290 278313
rect 123656 278161 124210 278177
rect 123656 278127 123672 278161
rect 124194 278127 124210 278161
rect 123656 278080 124210 278127
rect 122414 277745 123290 277792
rect 122414 277711 122430 277745
rect 123274 277711 123290 277745
rect 122414 277695 123290 277711
rect 122416 277581 123216 277597
rect 122416 277547 122432 277581
rect 123200 277547 123216 277581
rect 122416 277500 123216 277547
rect 122416 277353 123216 277400
rect 122416 277319 122432 277353
rect 123200 277319 123216 277353
rect 122416 277303 123216 277319
rect 123656 277347 124210 277394
rect 123656 277313 123672 277347
rect 124194 277313 124210 277347
rect 123656 277297 124210 277313
rect 122438 276749 123832 276765
rect 122438 276715 122454 276749
rect 123816 276715 123832 276749
rect 122438 276668 123832 276715
rect 122438 276445 123832 276492
rect 122438 276411 122454 276445
rect 123816 276411 123832 276445
rect 122438 276395 123832 276411
rect 122369 275795 122466 275811
rect 122369 275727 122385 275795
rect 122419 275727 122466 275795
rect 122369 275711 122466 275727
rect 122866 275795 122963 275811
rect 122866 275727 122913 275795
rect 122947 275727 122963 275795
rect 122866 275711 122963 275727
rect 123005 275795 123102 275811
rect 123005 275727 123021 275795
rect 123055 275727 123102 275795
rect 123005 275711 123102 275727
rect 123502 275795 123599 275811
rect 123502 275727 123549 275795
rect 123583 275727 123599 275795
rect 123502 275711 123599 275727
rect 123641 275795 123738 275811
rect 123641 275727 123657 275795
rect 123691 275727 123738 275795
rect 123641 275711 123738 275727
rect 124138 275795 124235 275811
rect 124138 275727 124185 275795
rect 124219 275727 124235 275795
rect 124138 275711 124235 275727
rect 124277 275795 124374 275811
rect 124277 275727 124293 275795
rect 124327 275727 124374 275795
rect 124277 275711 124374 275727
rect 124774 275795 124871 275811
rect 124774 275727 124821 275795
rect 124855 275727 124871 275795
rect 124774 275711 124871 275727
rect 122952 274934 123952 274950
rect 122952 274900 122968 274934
rect 123936 274900 123952 274934
rect 122952 274862 123952 274900
rect 122952 274624 123952 274662
rect 122952 274590 122968 274624
rect 123936 274590 123952 274624
rect 122952 274574 123952 274590
rect 122277 274350 122477 274366
rect 122277 274316 122293 274350
rect 122461 274316 122477 274350
rect 122277 274278 122477 274316
rect 122693 274350 122893 274366
rect 122693 274316 122709 274350
rect 122877 274316 122893 274350
rect 122693 274278 122893 274316
rect 123109 274350 123309 274366
rect 123109 274316 123125 274350
rect 123293 274316 123309 274350
rect 123109 274278 123309 274316
rect 123525 274350 123725 274366
rect 123525 274316 123541 274350
rect 123709 274316 123725 274350
rect 123525 274278 123725 274316
rect 123941 274350 124141 274366
rect 123941 274316 123957 274350
rect 124125 274316 124141 274350
rect 123941 274278 124141 274316
rect 124357 274350 124557 274366
rect 124357 274316 124373 274350
rect 124541 274316 124557 274350
rect 124357 274278 124557 274316
rect 122277 273740 122477 273778
rect 122277 273706 122293 273740
rect 122461 273706 122477 273740
rect 122277 273690 122477 273706
rect 122693 273740 122893 273778
rect 122693 273706 122709 273740
rect 122877 273706 122893 273740
rect 122693 273690 122893 273706
rect 123109 273740 123309 273778
rect 123109 273706 123125 273740
rect 123293 273706 123309 273740
rect 123109 273690 123309 273706
rect 123525 273740 123725 273778
rect 123525 273706 123541 273740
rect 123709 273706 123725 273740
rect 123525 273690 123725 273706
rect 123941 273740 124141 273778
rect 123941 273706 123957 273740
rect 124125 273706 124141 273740
rect 123941 273690 124141 273706
rect 124357 273740 124557 273778
rect 124357 273706 124373 273740
rect 124541 273706 124557 273740
rect 124357 273690 124557 273706
rect 122125 272894 122525 272910
rect 122125 272860 122141 272894
rect 122509 272860 122525 272894
rect 122125 272813 122525 272860
rect 122825 272894 123225 272910
rect 122825 272860 122841 272894
rect 123209 272860 123225 272894
rect 122825 272813 123225 272860
rect 122125 272666 122525 272713
rect 122125 272632 122141 272666
rect 122509 272632 122525 272666
rect 122125 272616 122525 272632
rect 122825 272666 123225 272713
rect 122825 272632 122841 272666
rect 123209 272632 123225 272666
rect 122825 272616 123225 272632
rect 122125 272510 122525 272526
rect 122125 272476 122141 272510
rect 122509 272476 122525 272510
rect 122125 272429 122525 272476
rect 122825 272510 123225 272526
rect 122825 272476 122841 272510
rect 123209 272476 123225 272510
rect 122825 272429 123225 272476
rect 122125 271882 122525 271929
rect 122125 271848 122141 271882
rect 122509 271848 122525 271882
rect 122125 271832 122525 271848
rect 122825 271882 123225 271929
rect 122825 271848 122841 271882
rect 123209 271848 123225 271882
rect 122825 271832 123225 271848
rect 122125 271726 122525 271742
rect 122125 271692 122141 271726
rect 122509 271692 122525 271726
rect 122125 271645 122525 271692
rect 122825 271726 123225 271742
rect 122825 271692 122841 271726
rect 123209 271692 123225 271726
rect 122825 271645 123225 271692
rect 122125 271098 122525 271145
rect 122125 271064 122141 271098
rect 122509 271064 122525 271098
rect 122125 271048 122525 271064
rect 122825 271098 123225 271145
rect 122825 271064 122841 271098
rect 123209 271064 123225 271098
rect 122825 271048 123225 271064
rect 122125 270942 122525 270958
rect 122125 270908 122141 270942
rect 122509 270908 122525 270942
rect 122125 270861 122525 270908
rect 122825 270942 123225 270958
rect 122825 270908 122841 270942
rect 123209 270908 123225 270942
rect 122825 270861 123225 270908
rect 122125 270314 122525 270361
rect 122125 270280 122141 270314
rect 122509 270280 122525 270314
rect 122125 270264 122525 270280
rect 122825 270314 123225 270361
rect 122825 270280 122841 270314
rect 123209 270280 123225 270314
rect 122825 270264 123225 270280
rect 122125 270158 122525 270174
rect 122125 270124 122141 270158
rect 122509 270124 122525 270158
rect 122125 270077 122525 270124
rect 122825 270158 123225 270174
rect 122825 270124 122841 270158
rect 123209 270124 123225 270158
rect 122825 270077 123225 270124
rect 122125 269530 122525 269577
rect 122125 269496 122141 269530
rect 122509 269496 122525 269530
rect 122125 269480 122525 269496
rect 122825 269530 123225 269577
rect 122825 269496 122841 269530
rect 123209 269496 123225 269530
rect 122825 269480 123225 269496
rect 122125 269374 122525 269390
rect 122125 269340 122141 269374
rect 122509 269340 122525 269374
rect 122125 269293 122525 269340
rect 122825 269374 123225 269390
rect 122825 269340 122841 269374
rect 123209 269340 123225 269374
rect 122825 269293 123225 269340
rect 122125 269146 122525 269193
rect 122125 269112 122141 269146
rect 122509 269112 122525 269146
rect 122125 269096 122525 269112
rect 122825 269146 123225 269193
rect 122825 269112 122841 269146
rect 123209 269112 123225 269146
rect 122825 269096 123225 269112
rect 124104 272504 124192 272520
rect 124104 272336 124120 272504
rect 124154 272336 124192 272504
rect 124104 272320 124192 272336
rect 124692 272504 124780 272520
rect 124692 272336 124730 272504
rect 124764 272336 124780 272504
rect 124692 272320 124780 272336
rect 124104 272088 124192 272104
rect 124104 271920 124120 272088
rect 124154 271920 124192 272088
rect 124104 271904 124192 271920
rect 124692 272088 124780 272104
rect 124692 271920 124730 272088
rect 124764 271920 124780 272088
rect 124692 271904 124780 271920
rect 124104 271672 124192 271688
rect 124104 271504 124120 271672
rect 124154 271504 124192 271672
rect 124104 271488 124192 271504
rect 124692 271672 124780 271688
rect 124692 271504 124730 271672
rect 124764 271504 124780 271672
rect 124692 271488 124780 271504
rect 124104 271256 124192 271272
rect 124104 271088 124120 271256
rect 124154 271088 124192 271256
rect 124104 271072 124192 271088
rect 124692 271256 124780 271272
rect 124692 271088 124730 271256
rect 124764 271088 124780 271256
rect 124692 271072 124780 271088
rect 124104 270840 124192 270856
rect 124104 270672 124120 270840
rect 124154 270672 124192 270840
rect 124104 270656 124192 270672
rect 124692 270840 124780 270856
rect 124692 270672 124730 270840
rect 124764 270672 124780 270840
rect 124692 270656 124780 270672
rect 124104 270424 124192 270440
rect 124104 270256 124120 270424
rect 124154 270256 124192 270424
rect 124104 270240 124192 270256
rect 124692 270424 124780 270440
rect 124692 270256 124730 270424
rect 124764 270256 124780 270424
rect 124692 270240 124780 270256
rect 124104 270008 124192 270024
rect 124104 269840 124120 270008
rect 124154 269840 124192 270008
rect 124104 269824 124192 269840
rect 124692 270008 124780 270024
rect 124692 269840 124730 270008
rect 124764 269840 124780 270008
rect 124692 269824 124780 269840
rect 124104 269592 124192 269608
rect 124104 269424 124120 269592
rect 124154 269424 124192 269592
rect 124104 269408 124192 269424
rect 124692 269592 124780 269608
rect 124692 269424 124730 269592
rect 124764 269424 124780 269592
rect 124692 269408 124780 269424
<< polycont >>
rect 106373 280851 106473 280885
rect 106773 280851 106873 280885
rect 107173 280851 107273 280885
rect 107573 280851 107673 280885
rect 107973 280851 108073 280885
rect 108373 280851 108473 280885
rect 108773 280851 108873 280885
rect 109173 280851 109273 280885
rect 109573 280851 109673 280885
rect 109973 280851 110073 280885
rect 106373 279721 106473 279755
rect 106773 279721 106873 279755
rect 107173 279721 107273 279755
rect 107573 279721 107673 279755
rect 107973 279721 108073 279755
rect 108373 279721 108473 279755
rect 108773 279721 108873 279755
rect 109173 279721 109273 279755
rect 109573 279721 109673 279755
rect 109973 279721 110073 279755
rect 106287 278773 106321 278995
rect 107629 278773 107663 278995
rect 106287 278173 106321 278395
rect 107629 278173 107663 278395
rect 106410 277106 106444 277148
rect 107572 277106 107606 277148
rect 109793 279049 110047 279083
rect 109793 277901 110047 277935
rect 109793 277793 110047 277827
rect 109793 276645 110047 276679
rect 106870 274951 106904 275697
rect 107176 274951 107210 275697
rect 107370 274951 107404 275697
rect 107676 274951 107710 275697
rect 107870 274951 107904 275697
rect 108176 274951 108210 275697
rect 108370 274951 108404 275697
rect 108676 274951 108710 275697
rect 108870 274951 108904 275697
rect 109176 274951 109210 275697
rect 109370 274951 109404 275697
rect 109676 274951 109710 275697
rect 107475 272117 108063 272151
rect 106997 272009 107175 272043
rect 106997 271735 107175 271769
rect 107475 271663 108063 271697
rect 107101 271327 107135 271473
rect 108411 271327 108445 271473
rect 107101 270957 107135 271103
rect 108411 270957 108445 271103
rect 109456 272473 109494 272507
rect 109456 270625 109494 270659
rect 111452 280676 111486 280804
rect 112662 280676 112696 280804
rect 112898 280644 112932 280812
rect 114108 280644 114142 280812
rect 111452 280316 111486 280444
rect 112662 280316 112696 280444
rect 112898 280220 112932 280388
rect 114108 280220 114142 280388
rect 111452 279956 111486 280084
rect 112662 279956 112696 280084
rect 112928 279938 112962 279986
rect 114138 279938 114172 279986
rect 111452 279596 111486 279724
rect 112662 279596 112696 279724
rect 112928 279640 112962 279688
rect 114138 279640 114172 279688
rect 114576 280419 114610 280787
rect 114904 280419 114938 280787
rect 114576 279973 114610 280101
rect 114904 279973 114938 280101
rect 114576 279565 114610 279693
rect 114904 279565 114938 279693
rect 115267 280419 115301 280787
rect 115595 280419 115629 280787
rect 115267 279973 115301 280101
rect 115595 279973 115629 280101
rect 115267 279565 115301 279693
rect 115595 279565 115629 279693
rect 116063 280644 116097 280812
rect 117273 280644 117307 280812
rect 117509 280676 117543 280804
rect 118719 280676 118753 280804
rect 116063 280220 116097 280388
rect 117273 280220 117307 280388
rect 117509 280316 117543 280444
rect 118719 280316 118753 280444
rect 116033 279938 116067 279986
rect 117243 279938 117277 279986
rect 117509 279956 117543 280084
rect 118719 279956 118753 280084
rect 116033 279640 116067 279688
rect 117243 279640 117277 279688
rect 117509 279596 117543 279724
rect 118719 279596 118753 279724
rect 111452 279010 111486 279138
rect 112662 279010 112696 279138
rect 112898 278978 112932 279146
rect 114108 278978 114142 279146
rect 111452 278650 111486 278778
rect 112662 278650 112696 278778
rect 112898 278554 112932 278722
rect 114108 278554 114142 278722
rect 111452 278290 111486 278418
rect 112662 278290 112696 278418
rect 112928 278272 112962 278320
rect 114138 278272 114172 278320
rect 111452 277930 111486 278058
rect 112662 277930 112696 278058
rect 112928 277974 112962 278022
rect 114138 277974 114172 278022
rect 114576 278753 114610 279121
rect 114904 278753 114938 279121
rect 114576 278307 114610 278435
rect 114904 278307 114938 278435
rect 114576 277899 114610 278027
rect 114904 277899 114938 278027
rect 115267 278753 115301 279121
rect 115595 278753 115629 279121
rect 115267 278307 115301 278435
rect 115595 278307 115629 278435
rect 115267 277899 115301 278027
rect 115595 277899 115629 278027
rect 116063 278978 116097 279146
rect 117273 278978 117307 279146
rect 117509 279010 117543 279138
rect 118719 279010 118753 279138
rect 116063 278554 116097 278722
rect 117273 278554 117307 278722
rect 117509 278650 117543 278778
rect 118719 278650 118753 278778
rect 116033 278272 116067 278320
rect 117243 278272 117277 278320
rect 117509 278290 117543 278418
rect 118719 278290 118753 278418
rect 116033 277974 116067 278022
rect 117243 277974 117277 278022
rect 117509 277930 117543 278058
rect 118719 277930 118753 278058
rect 111452 277344 111486 277472
rect 112662 277344 112696 277472
rect 112898 277312 112932 277480
rect 114108 277312 114142 277480
rect 111452 276984 111486 277112
rect 112662 276984 112696 277112
rect 112898 276888 112932 277056
rect 114108 276888 114142 277056
rect 111452 276624 111486 276752
rect 112662 276624 112696 276752
rect 112928 276606 112962 276654
rect 114138 276606 114172 276654
rect 111452 276264 111486 276392
rect 112662 276264 112696 276392
rect 112928 276308 112962 276356
rect 114138 276308 114172 276356
rect 114576 277087 114610 277455
rect 114904 277087 114938 277455
rect 114576 276641 114610 276769
rect 114904 276641 114938 276769
rect 114576 276233 114610 276361
rect 114904 276233 114938 276361
rect 115267 277087 115301 277455
rect 115595 277087 115629 277455
rect 115267 276641 115301 276769
rect 115595 276641 115629 276769
rect 115267 276233 115301 276361
rect 115595 276233 115629 276361
rect 116063 277312 116097 277480
rect 117273 277312 117307 277480
rect 117509 277344 117543 277472
rect 118719 277344 118753 277472
rect 116063 276888 116097 277056
rect 117273 276888 117307 277056
rect 117509 276984 117543 277112
rect 118719 276984 118753 277112
rect 116033 276606 116067 276654
rect 117243 276606 117277 276654
rect 117509 276624 117543 276752
rect 118719 276624 118753 276752
rect 116033 276308 116067 276356
rect 117243 276308 117277 276356
rect 117509 276264 117543 276392
rect 118719 276264 118753 276392
rect 111452 275678 111486 275806
rect 112662 275678 112696 275806
rect 112898 275646 112932 275814
rect 114108 275646 114142 275814
rect 111452 275318 111486 275446
rect 112662 275318 112696 275446
rect 112898 275222 112932 275390
rect 114108 275222 114142 275390
rect 111452 274958 111486 275086
rect 112662 274958 112696 275086
rect 112928 274940 112962 274988
rect 114138 274940 114172 274988
rect 111452 274598 111486 274726
rect 112662 274598 112696 274726
rect 112928 274642 112962 274690
rect 114138 274642 114172 274690
rect 114576 275421 114610 275789
rect 114904 275421 114938 275789
rect 114576 274975 114610 275103
rect 114904 274975 114938 275103
rect 114576 274567 114610 274695
rect 114904 274567 114938 274695
rect 115267 275421 115301 275789
rect 115595 275421 115629 275789
rect 115267 274975 115301 275103
rect 115595 274975 115629 275103
rect 115267 274567 115301 274695
rect 115595 274567 115629 274695
rect 116063 275646 116097 275814
rect 117273 275646 117307 275814
rect 117509 275678 117543 275806
rect 118719 275678 118753 275806
rect 116063 275222 116097 275390
rect 117273 275222 117307 275390
rect 117509 275318 117543 275446
rect 118719 275318 118753 275446
rect 116033 274940 116067 274988
rect 117243 274940 117277 274988
rect 117509 274958 117543 275086
rect 118719 274958 118753 275086
rect 116033 274642 116067 274690
rect 117243 274642 117277 274690
rect 117509 274598 117543 274726
rect 118719 274598 118753 274726
rect 111452 274012 111486 274140
rect 112662 274012 112696 274140
rect 112898 273980 112932 274148
rect 114108 273980 114142 274148
rect 111452 273652 111486 273780
rect 112662 273652 112696 273780
rect 112898 273556 112932 273724
rect 114108 273556 114142 273724
rect 111452 273292 111486 273420
rect 112662 273292 112696 273420
rect 112928 273274 112962 273322
rect 114138 273274 114172 273322
rect 111452 272932 111486 273060
rect 112662 272932 112696 273060
rect 112928 272976 112962 273024
rect 114138 272976 114172 273024
rect 114576 273755 114610 274123
rect 114904 273755 114938 274123
rect 114576 273309 114610 273437
rect 114904 273309 114938 273437
rect 114576 272901 114610 273029
rect 114904 272901 114938 273029
rect 115267 273755 115301 274123
rect 115595 273755 115629 274123
rect 115267 273309 115301 273437
rect 115595 273309 115629 273437
rect 115267 272901 115301 273029
rect 115595 272901 115629 273029
rect 116063 273980 116097 274148
rect 117273 273980 117307 274148
rect 117509 274012 117543 274140
rect 118719 274012 118753 274140
rect 116063 273556 116097 273724
rect 117273 273556 117307 273724
rect 117509 273652 117543 273780
rect 118719 273652 118753 273780
rect 116033 273274 116067 273322
rect 117243 273274 117277 273322
rect 117509 273292 117543 273420
rect 118719 273292 118753 273420
rect 116033 272976 116067 273024
rect 117243 272976 117277 273024
rect 117509 272932 117543 273060
rect 118719 272932 118753 273060
rect 115897 271962 116025 271996
rect 116297 271962 116425 271996
rect 116697 271962 116825 271996
rect 117097 271962 117225 271996
rect 117497 271962 117625 271996
rect 117897 271962 118025 271996
rect 118297 271962 118425 271996
rect 118697 271962 118825 271996
rect 112594 271353 112722 271387
rect 112994 271353 113122 271387
rect 113394 271353 113522 271387
rect 113794 271353 113922 271387
rect 112594 271025 112722 271059
rect 112994 271025 113122 271059
rect 113394 271025 113522 271059
rect 113794 271025 113922 271059
rect 114653 271324 114781 271358
rect 115053 271324 115181 271358
rect 114653 270996 114781 271030
rect 115053 270996 115181 271030
rect 115897 270752 116025 270786
rect 116297 270752 116425 270786
rect 116697 270752 116825 270786
rect 117097 270752 117225 270786
rect 117497 270752 117625 270786
rect 117897 270752 118025 270786
rect 118297 270752 118425 270786
rect 118697 270752 118825 270786
rect 112576 270262 112704 270296
rect 112976 270262 113104 270296
rect 113376 270262 113504 270296
rect 113776 270262 113904 270296
rect 114176 270262 114304 270296
rect 114576 270262 114704 270296
rect 114976 270262 115104 270296
rect 115376 270262 115504 270296
rect 115776 270262 115904 270296
rect 116176 270262 116304 270296
rect 116576 270262 116704 270296
rect 116976 270262 117104 270296
rect 117376 270262 117504 270296
rect 117776 270262 117904 270296
rect 118176 270262 118304 270296
rect 118576 270262 118704 270296
rect 112576 269052 112704 269086
rect 112976 269052 113104 269086
rect 113376 269052 113504 269086
rect 113776 269052 113904 269086
rect 114176 269052 114304 269086
rect 114576 269052 114704 269086
rect 114976 269052 115104 269086
rect 115376 269052 115504 269086
rect 115776 269052 115904 269086
rect 116176 269052 116304 269086
rect 116576 269052 116704 269086
rect 116976 269052 117104 269086
rect 117376 269052 117504 269086
rect 117776 269052 117904 269086
rect 118176 269052 118304 269086
rect 118576 269052 118704 269086
rect 120445 280684 120813 280718
rect 121145 280684 121513 280718
rect 120445 280456 120813 280490
rect 121145 280456 121513 280490
rect 120445 280300 120813 280334
rect 121145 280300 121513 280334
rect 120445 279672 120813 279706
rect 121145 279672 121513 279706
rect 120445 279516 120813 279550
rect 121145 279516 121513 279550
rect 120445 278888 120813 278922
rect 121145 278888 121513 278922
rect 120445 278732 120813 278766
rect 121145 278732 121513 278766
rect 120445 278104 120813 278138
rect 121145 278104 121513 278138
rect 120445 277948 120813 277982
rect 121145 277948 121513 277982
rect 120445 277320 120813 277354
rect 121145 277320 121513 277354
rect 120445 277164 120813 277198
rect 121145 277164 121513 277198
rect 120445 276536 120813 276570
rect 121145 276536 121513 276570
rect 120445 276380 120813 276414
rect 121145 276380 121513 276414
rect 120445 275752 120813 275786
rect 121145 275752 121513 275786
rect 120445 275596 120813 275630
rect 121145 275596 121513 275630
rect 120445 274968 120813 275002
rect 121145 274968 121513 275002
rect 120445 274812 120813 274846
rect 121145 274812 121513 274846
rect 120445 274184 120813 274218
rect 121145 274184 121513 274218
rect 120445 274028 120813 274062
rect 121145 274028 121513 274062
rect 120445 273400 120813 273434
rect 121145 273400 121513 273434
rect 120445 273244 120813 273278
rect 121145 273244 121513 273278
rect 120445 272616 120813 272650
rect 121145 272616 121513 272650
rect 120445 272460 120813 272494
rect 121145 272460 121513 272494
rect 120445 271832 120813 271866
rect 121145 271832 121513 271866
rect 120445 271676 120813 271710
rect 121145 271676 121513 271710
rect 120445 271048 120813 271082
rect 121145 271048 121513 271082
rect 120445 270892 120813 270926
rect 121145 270892 121513 270926
rect 120445 270264 120813 270298
rect 121145 270264 121513 270298
rect 120445 270108 120813 270142
rect 121145 270108 121513 270142
rect 120445 269480 120813 269514
rect 121145 269480 121513 269514
rect 120445 269324 120813 269358
rect 121145 269324 121513 269358
rect 120445 269096 120813 269130
rect 121145 269096 121513 269130
rect 122372 280470 122740 280504
rect 123072 280470 123440 280504
rect 122372 279842 122740 279876
rect 123072 279842 123440 279876
rect 122372 279686 122740 279720
rect 123072 279686 123440 279720
rect 122372 279058 122740 279092
rect 123072 279058 123440 279092
rect 122430 278313 123274 278347
rect 123672 278127 124194 278161
rect 122430 277711 123274 277745
rect 122432 277547 123200 277581
rect 122432 277319 123200 277353
rect 123672 277313 124194 277347
rect 122454 276715 123816 276749
rect 122454 276411 123816 276445
rect 122385 275727 122419 275795
rect 122913 275727 122947 275795
rect 123021 275727 123055 275795
rect 123549 275727 123583 275795
rect 123657 275727 123691 275795
rect 124185 275727 124219 275795
rect 124293 275727 124327 275795
rect 124821 275727 124855 275795
rect 122968 274900 123936 274934
rect 122968 274590 123936 274624
rect 122293 274316 122461 274350
rect 122709 274316 122877 274350
rect 123125 274316 123293 274350
rect 123541 274316 123709 274350
rect 123957 274316 124125 274350
rect 124373 274316 124541 274350
rect 122293 273706 122461 273740
rect 122709 273706 122877 273740
rect 123125 273706 123293 273740
rect 123541 273706 123709 273740
rect 123957 273706 124125 273740
rect 124373 273706 124541 273740
rect 122141 272860 122509 272894
rect 122841 272860 123209 272894
rect 122141 272632 122509 272666
rect 122841 272632 123209 272666
rect 122141 272476 122509 272510
rect 122841 272476 123209 272510
rect 122141 271848 122509 271882
rect 122841 271848 123209 271882
rect 122141 271692 122509 271726
rect 122841 271692 123209 271726
rect 122141 271064 122509 271098
rect 122841 271064 123209 271098
rect 122141 270908 122509 270942
rect 122841 270908 123209 270942
rect 122141 270280 122509 270314
rect 122841 270280 123209 270314
rect 122141 270124 122509 270158
rect 122841 270124 123209 270158
rect 122141 269496 122509 269530
rect 122841 269496 123209 269530
rect 122141 269340 122509 269374
rect 122841 269340 123209 269374
rect 122141 269112 122509 269146
rect 122841 269112 123209 269146
rect 124120 272336 124154 272504
rect 124730 272336 124764 272504
rect 124120 271920 124154 272088
rect 124730 271920 124764 272088
rect 124120 271504 124154 271672
rect 124730 271504 124764 271672
rect 124120 271088 124154 271256
rect 124730 271088 124764 271256
rect 124120 270672 124154 270840
rect 124730 270672 124764 270840
rect 124120 270256 124154 270424
rect 124730 270256 124764 270424
rect 124120 269840 124154 270008
rect 124730 269840 124764 270008
rect 124120 269424 124154 269592
rect 124730 269424 124764 269592
<< locali >>
rect 125105 281915 125658 281925
rect 105823 281315 125658 281915
rect 105976 281064 106456 281315
rect 105974 281045 106456 281064
rect 108743 281045 110315 281315
rect 111807 281179 118652 281315
rect 105974 281041 106170 281045
rect 106060 280961 106170 281041
rect 110228 281005 110315 281045
rect 111046 281107 111234 281179
rect 110228 280961 110313 281005
rect 106060 280885 106465 280961
rect 106060 280880 106373 280885
rect 106060 279716 106125 280880
rect 106207 280851 106373 280880
rect 106473 280851 106489 280885
rect 106207 280801 106345 280851
rect 106666 280817 106711 280961
rect 106757 280851 106773 280885
rect 106873 280851 106889 280885
rect 107066 280817 107111 280961
rect 107157 280851 107173 280885
rect 107273 280851 107289 280885
rect 107466 280817 107511 280961
rect 107557 280851 107573 280885
rect 107673 280851 107689 280885
rect 107866 280817 107911 280961
rect 107957 280851 107973 280885
rect 108073 280851 108089 280885
rect 108357 280851 108373 280885
rect 108473 280851 108489 280885
rect 108535 280817 108580 280961
rect 108757 280851 108773 280885
rect 108873 280851 108889 280885
rect 108935 280817 108980 280961
rect 109157 280851 109173 280885
rect 109273 280851 109289 280885
rect 109335 280817 109380 280961
rect 109557 280851 109573 280885
rect 109673 280851 109689 280885
rect 109735 280817 109780 280961
rect 109980 280885 110313 280961
rect 109957 280851 109973 280885
rect 110073 280862 110313 280885
rect 110073 280851 110231 280862
rect 110129 280817 110231 280851
rect 106207 279805 106311 280801
rect 106207 279789 106345 279805
rect 106501 280801 106535 280817
rect 106501 279789 106535 279805
rect 106666 280801 106745 280817
rect 106666 279805 106711 280801
rect 106666 279789 106745 279805
rect 106901 280801 106935 280817
rect 106901 279789 106935 279805
rect 107066 280801 107145 280817
rect 107066 279805 107111 280801
rect 107066 279789 107145 279805
rect 107301 280801 107335 280817
rect 107301 279789 107335 279805
rect 107466 280801 107545 280817
rect 107466 279805 107511 280801
rect 107466 279789 107545 279805
rect 107701 280801 107735 280817
rect 107701 279789 107735 279805
rect 107866 280801 107945 280817
rect 107866 279805 107911 280801
rect 107866 279789 107945 279805
rect 108101 280801 108135 280817
rect 108101 279789 108135 279805
rect 108311 280801 108345 280817
rect 108311 279789 108345 279805
rect 108501 280801 108580 280817
rect 108535 279805 108580 280801
rect 108501 279789 108580 279805
rect 108711 280801 108745 280817
rect 108711 279789 108745 279805
rect 108901 280801 108980 280817
rect 108935 279805 108980 280801
rect 108901 279789 108980 279805
rect 109111 280801 109145 280817
rect 109111 279789 109145 279805
rect 109301 280801 109380 280817
rect 109335 279805 109380 280801
rect 109301 279789 109380 279805
rect 109511 280801 109545 280817
rect 109511 279789 109545 279805
rect 109701 280801 109780 280817
rect 109735 279805 109780 280801
rect 109701 279789 109780 279805
rect 109911 280801 109945 280817
rect 109911 279789 109945 279805
rect 110101 280801 110231 280817
rect 110135 279805 110231 280801
rect 110101 279789 110231 279805
rect 106207 279755 106326 279789
rect 106489 279755 106535 279789
rect 109911 279755 109957 279789
rect 106207 279721 106373 279755
rect 106473 279721 106535 279755
rect 106757 279721 106773 279755
rect 106873 279721 106889 279755
rect 107157 279721 107173 279755
rect 107273 279721 107289 279755
rect 107557 279721 107573 279755
rect 107673 279721 107689 279755
rect 107957 279721 107973 279755
rect 108073 279721 108089 279755
rect 108357 279721 108373 279755
rect 108473 279721 108489 279755
rect 108757 279721 108773 279755
rect 108873 279721 108889 279755
rect 109157 279721 109173 279755
rect 109273 279721 109289 279755
rect 109557 279721 109573 279755
rect 109673 279721 109689 279755
rect 109911 279721 109973 279755
rect 110073 279747 110089 279755
rect 110129 279747 110231 279789
rect 110073 279721 110231 279747
rect 106207 279716 106463 279721
rect 106060 279625 106463 279716
rect 106757 279687 109689 279721
rect 109982 279698 110231 279721
rect 109982 279625 110313 279698
rect 106060 279549 106170 279625
rect 106125 279541 106170 279549
rect 110228 279541 110313 279625
rect 106169 279188 106229 279222
rect 107708 279188 107768 279222
rect 106169 279162 106203 279188
rect 107734 279162 107768 279188
rect 109636 279185 110312 279541
rect 106364 279023 106380 279057
rect 107570 279023 107586 279057
rect 106275 278995 106321 279011
rect 106275 278773 106287 278995
rect 106275 278395 106321 278773
rect 107629 278995 107675 279011
rect 107663 278773 107675 278995
rect 106364 278711 106380 278745
rect 107570 278711 107586 278745
rect 106364 278423 106380 278457
rect 107570 278423 107586 278457
rect 106275 278173 106287 278395
rect 106275 278157 106321 278173
rect 107629 278395 107675 278773
rect 107663 278173 107675 278395
rect 107629 278157 107675 278173
rect 106364 278111 106380 278145
rect 107570 278111 107586 278145
rect 106169 277984 106203 278010
rect 106762 278068 107237 278111
rect 106762 277984 106941 278068
rect 107098 277984 107237 278068
rect 107734 277984 107768 278010
rect 106169 277950 106229 277984
rect 107708 277950 107768 277984
rect 109617 279151 109713 279185
rect 110127 279151 110312 279185
rect 109617 279089 109651 279151
rect 106902 277789 106941 277950
rect 107098 277789 107130 277950
rect 106902 277724 107130 277789
rect 106308 277290 106404 277324
rect 107612 277290 107708 277324
rect 106308 277228 106342 277290
rect 107674 277228 107708 277290
rect 106487 277176 106503 277210
rect 107513 277176 107529 277210
rect 106410 277148 106444 277164
rect 106410 277090 106444 277106
rect 107572 277148 107606 277164
rect 107572 277090 107606 277106
rect 106487 277044 106503 277078
rect 107513 277044 107529 277078
rect 106308 276964 106342 277026
rect 106849 276964 107133 277044
rect 107674 276964 107708 277026
rect 106308 276930 106404 276964
rect 107612 276930 107708 276964
rect 106719 276403 106985 276930
rect 110189 279089 110312 279151
rect 109777 279049 109793 279083
rect 110047 279049 110063 279083
rect 109731 278999 109765 279015
rect 109731 277969 109765 277985
rect 110075 278999 110109 279015
rect 110075 277969 110109 277985
rect 109777 277901 109793 277935
rect 110047 277901 110063 277935
rect 109777 277793 109793 277827
rect 110047 277793 110063 277827
rect 109731 277743 109765 277759
rect 109731 276713 109765 276729
rect 110075 277743 110109 277759
rect 110075 276713 110109 276729
rect 109777 276645 109793 276679
rect 110047 276645 110063 276679
rect 109617 276577 109651 276639
rect 110223 276639 110312 279089
rect 110189 276577 110312 276639
rect 109617 276543 109713 276577
rect 110127 276553 110312 276577
rect 110127 276543 110224 276553
rect 106294 276290 106985 276403
rect 106294 274853 106375 276290
rect 106549 275934 106985 276290
rect 110145 276056 110224 276543
rect 106549 275900 106766 275934
rect 109787 275900 109847 275934
rect 106549 275874 106887 275900
rect 106549 274853 106706 275874
rect 106294 274773 106706 274853
rect 106740 275713 106887 275874
rect 106995 275759 107075 275900
rect 109498 275759 109578 275900
rect 109693 275874 109847 275900
rect 106947 275725 106963 275759
rect 107117 275725 107133 275759
rect 107447 275725 107463 275759
rect 107617 275725 107633 275759
rect 107947 275725 107963 275759
rect 108117 275725 108133 275759
rect 108447 275725 108463 275759
rect 108617 275725 108633 275759
rect 108947 275725 108963 275759
rect 109117 275725 109133 275759
rect 109447 275725 109463 275759
rect 109617 275725 109633 275759
rect 109693 275713 109813 275874
rect 106740 275697 106904 275713
rect 106740 274951 106870 275697
rect 106740 274935 106904 274951
rect 107176 275697 107210 275713
rect 107176 274935 107210 274951
rect 107370 275697 107404 275713
rect 107370 274935 107404 274951
rect 107676 275697 107710 275713
rect 107676 274935 107710 274951
rect 107870 275697 107904 275713
rect 107870 274935 107904 274951
rect 108176 275697 108210 275713
rect 108176 274935 108210 274951
rect 108370 275697 108404 275713
rect 108370 274935 108404 274951
rect 108676 275697 108710 275713
rect 108676 274935 108710 274951
rect 108870 275697 108904 275713
rect 108870 274935 108904 274951
rect 109176 275697 109210 275713
rect 109176 274935 109210 274951
rect 109370 275697 109404 275713
rect 109370 274935 109404 274951
rect 109676 275697 109813 275713
rect 109710 274951 109813 275697
rect 109676 274935 109813 274951
rect 106740 274886 106891 274935
rect 106947 274889 106963 274923
rect 107117 274889 107133 274923
rect 107447 274889 107463 274923
rect 107617 274889 107633 274923
rect 107947 274889 107963 274923
rect 108117 274889 108133 274923
rect 108447 274889 108463 274923
rect 108617 274889 108633 274923
rect 108947 274889 108963 274923
rect 109117 274889 109133 274923
rect 109447 274889 109463 274923
rect 109617 274889 109633 274923
rect 106947 274886 109633 274889
rect 106740 274882 109633 274886
rect 109692 274882 109813 274935
rect 106740 274773 109813 274882
rect 106294 274747 109847 274773
rect 106294 274731 106766 274747
rect 106706 274713 106766 274731
rect 109787 274713 109847 274747
rect 105974 274619 106060 274635
rect 110145 274619 110224 274669
rect 105974 274527 106114 274619
rect 110167 274527 110224 274619
rect 106281 272918 106580 272951
rect 106459 272794 106580 272918
rect 109977 272918 110259 272951
rect 109977 272794 110081 272918
rect 106459 272786 110081 272794
rect 107343 272367 108250 272786
rect 109088 272568 109148 272602
rect 109801 272568 109861 272602
rect 109088 272542 109122 272568
rect 106715 272339 106843 272367
rect 106789 272299 106843 272339
rect 106887 272299 106963 272367
rect 108657 272339 108803 272367
rect 108657 272299 108729 272339
rect 107459 272117 107475 272151
rect 108063 272117 108079 272151
rect 107413 272067 107447 272083
rect 106981 272009 106997 272043
rect 107175 272009 107191 272043
rect 106789 271959 106969 271975
rect 106789 271819 106935 271959
rect 106789 271803 106969 271819
rect 107203 271959 107237 271975
rect 107203 271803 107237 271819
rect 106981 271735 106997 271769
rect 107175 271735 107191 271769
rect 107413 271731 107447 271747
rect 108091 272067 108125 272083
rect 108091 271731 108125 271747
rect 107459 271663 107475 271697
rect 108063 271663 108079 271697
rect 107169 271501 107185 271535
rect 108361 271501 108377 271535
rect 107101 271473 107135 271489
rect 107101 271311 107135 271327
rect 108411 271473 108445 271489
rect 108411 271311 108445 271327
rect 107169 271265 107185 271299
rect 108361 271265 108377 271299
rect 107169 271131 107185 271165
rect 108361 271131 108377 271165
rect 107101 271103 107135 271119
rect 107101 270941 107135 270957
rect 108411 271103 108445 271119
rect 108411 270941 108445 270957
rect 107169 270895 107185 270929
rect 108361 270895 108377 270929
rect 106789 270773 106869 270801
rect 106715 270733 106869 270773
rect 108683 270773 108729 270801
rect 108947 271005 109088 271029
rect 108947 270837 108976 271005
rect 109077 270837 109088 271005
rect 108947 270811 109088 270837
rect 108683 270733 108803 270773
rect 107329 270334 108364 270733
rect 109827 272542 109861 272568
rect 109394 272473 109456 272507
rect 109494 272473 109556 272507
rect 109394 272414 109428 272473
rect 109394 270659 109428 270718
rect 109522 272414 109556 272473
rect 109522 270659 109556 270718
rect 109394 270625 109456 270659
rect 109494 270625 109556 270659
rect 109088 270555 109122 270581
rect 109827 270555 109861 270581
rect 109088 270521 109148 270555
rect 109801 270521 109861 270555
rect 106459 270193 106570 270334
rect 106281 270177 106570 270193
rect 109967 270193 110081 270334
rect 111200 281099 111234 281107
rect 118876 281107 119159 281179
rect 122520 281165 125658 281315
rect 118876 281099 119005 281107
rect 113036 280904 114022 281099
rect 114455 280929 114515 280963
rect 115001 280929 115204 280963
rect 115690 280929 115750 280963
rect 111520 280866 112814 280902
rect 113036 280900 114246 280904
rect 114455 280903 114489 280929
rect 113036 280899 114353 280900
rect 111520 280832 111536 280866
rect 112612 280832 112628 280866
rect 111452 280804 111486 280820
rect 111452 280660 111486 280676
rect 112662 280804 112696 280820
rect 112662 280660 112696 280676
rect 111520 280614 111536 280648
rect 112612 280614 112628 280648
rect 111334 280578 112628 280614
rect 112772 280582 112814 280866
rect 112966 280884 114353 280899
rect 112966 280874 114235 280884
rect 112966 280840 112982 280874
rect 114058 280870 114235 280874
rect 114058 280840 114074 280870
rect 112898 280812 112932 280828
rect 112898 280628 112932 280644
rect 114108 280812 114142 280828
rect 114108 280628 114142 280644
rect 114210 280766 114235 280870
rect 114210 280750 114353 280766
rect 112966 280582 112982 280616
rect 114058 280582 114074 280616
rect 111334 280254 111376 280578
rect 112772 280548 114074 280582
rect 112772 280542 112832 280548
rect 111520 280506 112832 280542
rect 111520 280472 111536 280506
rect 112612 280472 112628 280506
rect 111452 280444 111486 280460
rect 111452 280300 111486 280316
rect 112662 280444 112696 280460
rect 112662 280300 112696 280316
rect 111520 280254 111536 280288
rect 112612 280254 112628 280288
rect 111334 280218 112628 280254
rect 111334 279894 111376 280218
rect 112772 280182 112832 280506
rect 114210 280484 114246 280750
rect 112966 280450 114246 280484
rect 112966 280416 112982 280450
rect 114058 280416 114074 280450
rect 112898 280388 112932 280404
rect 112898 280204 112932 280220
rect 114108 280388 114142 280404
rect 114108 280204 114142 280220
rect 111520 280160 112832 280182
rect 112966 280160 112982 280192
rect 111520 280158 112982 280160
rect 114058 280158 114074 280192
rect 111520 280146 114074 280158
rect 111520 280112 111536 280146
rect 112612 280112 112628 280146
rect 112744 280143 114074 280146
rect 112744 280126 114396 280143
rect 111452 280084 111486 280100
rect 111452 279940 111486 279956
rect 112662 280084 112696 280100
rect 112662 279940 112696 279956
rect 111520 279894 111536 279928
rect 112612 279894 112628 279928
rect 111334 279858 112628 279894
rect 111334 279534 111376 279858
rect 112744 279822 112780 280126
rect 113892 280107 114396 280126
rect 111520 279786 112780 279822
rect 112832 280048 113264 280082
rect 112832 280040 113012 280048
rect 112832 279786 112872 280040
rect 112996 280014 113012 280040
rect 114088 280014 114104 280048
rect 112928 279986 112962 280002
rect 112928 279922 112962 279938
rect 114138 279986 114172 280002
rect 114138 279922 114172 279938
rect 114324 279976 114396 280107
rect 112996 279882 113012 279910
rect 112994 279876 113012 279882
rect 114088 279882 114104 279910
rect 114324 279893 114342 279976
rect 114377 279893 114396 279976
rect 114088 279876 114274 279882
rect 112994 279836 114274 279876
rect 114324 279869 114396 279893
rect 111520 279752 111536 279786
rect 112612 279752 112628 279786
rect 112832 279750 113216 279786
rect 112832 279746 113012 279750
rect 111452 279724 111486 279740
rect 111452 279580 111486 279596
rect 112662 279724 112696 279740
rect 112832 279718 112872 279746
rect 112996 279716 113012 279746
rect 114088 279716 114104 279750
rect 112928 279688 112962 279704
rect 112928 279624 112962 279640
rect 114138 279688 114172 279704
rect 114138 279624 114172 279640
rect 112662 279580 112696 279596
rect 112996 279578 113012 279612
rect 114088 279578 114104 279612
rect 114234 279578 114274 279836
rect 111520 279534 111536 279568
rect 112612 279534 112628 279568
rect 111334 279498 112628 279534
rect 112994 279532 114455 279578
rect 113982 279425 114266 279430
rect 111312 279335 111328 279425
rect 114242 279335 114266 279425
rect 114652 280849 114862 280929
rect 114652 280815 114669 280849
rect 114845 280815 114862 280849
rect 114652 280814 114862 280815
rect 115027 280903 115178 280929
rect 114576 280787 114610 280803
rect 114576 280275 114610 280419
rect 114904 280787 114938 280803
rect 114653 280357 114669 280391
rect 114845 280357 114861 280391
rect 114904 280311 114938 280419
rect 114865 280294 114970 280311
rect 114865 280275 114885 280294
rect 114576 280227 114885 280275
rect 114576 280101 114610 280227
rect 114865 280226 114885 280227
rect 114948 280226 114970 280294
rect 114865 280204 114970 280226
rect 114653 280129 114669 280163
rect 114845 280129 114861 280163
rect 114576 279957 114610 279973
rect 114904 280101 114938 280204
rect 114904 279957 114938 279973
rect 114653 279911 114669 279945
rect 114845 279911 114861 279945
rect 114653 279874 114709 279911
rect 114805 279876 114861 279911
rect 114538 279835 114709 279874
rect 114804 279861 114991 279876
rect 114538 279709 114576 279835
rect 114804 279813 114868 279861
rect 114965 279813 114991 279861
rect 114804 279791 114991 279813
rect 114653 279721 114669 279755
rect 114845 279721 114861 279755
rect 114938 279709 114975 279791
rect 114538 279693 114610 279709
rect 114538 279565 114576 279693
rect 114538 279549 114610 279565
rect 114904 279693 114975 279709
rect 114938 279565 114975 279693
rect 114904 279549 114975 279565
rect 114653 279503 114669 279537
rect 114845 279503 114861 279537
rect 114455 279403 114489 279429
rect 114930 279429 115027 279487
rect 115061 279429 115144 280903
rect 115343 280849 115553 280929
rect 115343 280815 115360 280849
rect 115536 280815 115553 280849
rect 115343 280814 115553 280815
rect 115716 280903 115750 280929
rect 116183 280904 117169 281099
rect 115267 280787 115301 280803
rect 115267 280311 115301 280419
rect 115595 280787 115629 280803
rect 115344 280357 115360 280391
rect 115536 280357 115552 280391
rect 115235 280294 115340 280311
rect 115235 280226 115257 280294
rect 115320 280275 115340 280294
rect 115595 280275 115629 280419
rect 115320 280227 115629 280275
rect 115320 280226 115340 280227
rect 115235 280204 115340 280226
rect 115267 280101 115301 280204
rect 115344 280129 115360 280163
rect 115536 280129 115552 280163
rect 115267 279957 115301 279973
rect 115595 280101 115629 280227
rect 115595 279957 115629 279973
rect 115344 279911 115360 279945
rect 115536 279911 115552 279945
rect 115344 279876 115400 279911
rect 115214 279861 115401 279876
rect 115214 279813 115240 279861
rect 115337 279813 115401 279861
rect 115496 279874 115552 279911
rect 115496 279835 115667 279874
rect 115214 279791 115401 279813
rect 115230 279709 115267 279791
rect 115344 279721 115360 279755
rect 115536 279721 115552 279755
rect 115629 279709 115667 279835
rect 115230 279693 115301 279709
rect 115230 279565 115267 279693
rect 115230 279549 115301 279565
rect 115595 279693 115667 279709
rect 115629 279565 115667 279693
rect 115595 279549 115667 279565
rect 115344 279503 115360 279537
rect 115536 279503 115552 279537
rect 115178 279429 115275 279487
rect 114930 279403 115275 279429
rect 115959 280900 117169 280904
rect 115852 280899 117169 280900
rect 115852 280884 117239 280899
rect 115970 280874 117239 280884
rect 115970 280870 116147 280874
rect 115970 280766 115995 280870
rect 116131 280840 116147 280870
rect 117223 280840 117239 280874
rect 117391 280866 118685 280902
rect 115852 280750 115995 280766
rect 115959 280484 115995 280750
rect 116063 280812 116097 280828
rect 116063 280628 116097 280644
rect 117273 280812 117307 280828
rect 117273 280628 117307 280644
rect 116131 280582 116147 280616
rect 117223 280582 117239 280616
rect 117391 280582 117433 280866
rect 117577 280832 117593 280866
rect 118669 280832 118685 280866
rect 117509 280804 117543 280820
rect 117509 280660 117543 280676
rect 118719 280804 118753 280820
rect 118719 280660 118753 280676
rect 116131 280548 117433 280582
rect 117577 280614 117593 280648
rect 118669 280614 118685 280648
rect 117577 280578 118871 280614
rect 117373 280542 117433 280548
rect 117373 280506 118685 280542
rect 115959 280450 117239 280484
rect 116131 280416 116147 280450
rect 117223 280416 117239 280450
rect 116063 280388 116097 280404
rect 116063 280204 116097 280220
rect 117273 280388 117307 280404
rect 117273 280204 117307 280220
rect 116131 280158 116147 280192
rect 117223 280160 117239 280192
rect 117373 280182 117433 280506
rect 117577 280472 117593 280506
rect 118669 280472 118685 280506
rect 117509 280444 117543 280460
rect 117509 280300 117543 280316
rect 118719 280444 118753 280460
rect 118719 280300 118753 280316
rect 117577 280254 117593 280288
rect 118669 280254 118685 280288
rect 118829 280254 118871 280578
rect 117577 280218 118871 280254
rect 117373 280160 118685 280182
rect 117223 280158 118685 280160
rect 116131 280146 118685 280158
rect 116131 280143 117461 280146
rect 115809 280126 117461 280143
rect 115809 280107 116313 280126
rect 115809 279976 115881 280107
rect 116941 280048 117373 280082
rect 116101 280014 116117 280048
rect 117193 280040 117373 280048
rect 117193 280014 117209 280040
rect 115809 279893 115828 279976
rect 115863 279893 115881 279976
rect 116033 279986 116067 280002
rect 116033 279922 116067 279938
rect 117243 279986 117277 280002
rect 117243 279922 117277 279938
rect 115809 279869 115881 279893
rect 116101 279882 116117 279910
rect 115931 279876 116117 279882
rect 117193 279882 117209 279910
rect 117193 279876 117211 279882
rect 115931 279836 117211 279876
rect 115931 279578 115971 279836
rect 117333 279786 117373 280040
rect 117425 279822 117461 280126
rect 117577 280112 117593 280146
rect 118669 280112 118685 280146
rect 117509 280084 117543 280100
rect 117509 279940 117543 279956
rect 118719 280084 118753 280100
rect 118719 279940 118753 279956
rect 117577 279894 117593 279928
rect 118669 279894 118685 279928
rect 118829 279894 118871 280218
rect 117577 279858 118871 279894
rect 117425 279786 118685 279822
rect 116989 279750 117373 279786
rect 117577 279752 117593 279786
rect 118669 279752 118685 279786
rect 116101 279716 116117 279750
rect 117193 279746 117373 279750
rect 117193 279716 117209 279746
rect 117333 279718 117373 279746
rect 117509 279724 117543 279740
rect 116033 279688 116067 279704
rect 116033 279624 116067 279640
rect 117243 279688 117277 279704
rect 117243 279624 117277 279640
rect 116101 279578 116117 279612
rect 117193 279578 117209 279612
rect 117509 279580 117543 279596
rect 118719 279724 118753 279740
rect 118719 279580 118753 279596
rect 115750 279532 117211 279578
rect 117577 279534 117593 279568
rect 118669 279534 118685 279568
rect 118829 279534 118871 279858
rect 117577 279498 118871 279534
rect 115716 279403 115750 279429
rect 114455 279369 114515 279403
rect 115001 279369 115204 279403
rect 115690 279369 115750 279403
rect 115939 279425 116223 279430
rect 113036 279330 114266 279335
rect 113036 279238 114022 279330
rect 115061 279297 115144 279369
rect 115939 279335 115963 279425
rect 118877 279335 118893 279425
rect 115939 279330 117169 279335
rect 114455 279263 114515 279297
rect 115001 279263 115204 279297
rect 115690 279263 115750 279297
rect 111520 279200 112814 279236
rect 113036 279234 114246 279238
rect 114455 279237 114489 279263
rect 113036 279233 114353 279234
rect 111520 279166 111536 279200
rect 112612 279166 112628 279200
rect 111452 279138 111486 279154
rect 111452 278994 111486 279010
rect 112662 279138 112696 279154
rect 112662 278994 112696 279010
rect 111520 278948 111536 278982
rect 112612 278948 112628 278982
rect 111334 278912 112628 278948
rect 112772 278916 112814 279200
rect 112966 279218 114353 279233
rect 112966 279208 114235 279218
rect 112966 279174 112982 279208
rect 114058 279204 114235 279208
rect 114058 279174 114074 279204
rect 112898 279146 112932 279162
rect 112898 278962 112932 278978
rect 114108 279146 114142 279162
rect 114108 278962 114142 278978
rect 114210 279100 114235 279204
rect 114210 279084 114353 279100
rect 112966 278916 112982 278950
rect 114058 278916 114074 278950
rect 111334 278588 111376 278912
rect 112772 278882 114074 278916
rect 112772 278876 112832 278882
rect 111520 278840 112832 278876
rect 111520 278806 111536 278840
rect 112612 278806 112628 278840
rect 111452 278778 111486 278794
rect 111452 278634 111486 278650
rect 112662 278778 112696 278794
rect 112662 278634 112696 278650
rect 111520 278588 111536 278622
rect 112612 278588 112628 278622
rect 111334 278552 112628 278588
rect 111334 278228 111376 278552
rect 112772 278516 112832 278840
rect 114210 278818 114246 279084
rect 112966 278784 114246 278818
rect 112966 278750 112982 278784
rect 114058 278750 114074 278784
rect 112898 278722 112932 278738
rect 112898 278538 112932 278554
rect 114108 278722 114142 278738
rect 114108 278538 114142 278554
rect 111520 278494 112832 278516
rect 112966 278494 112982 278526
rect 111520 278492 112982 278494
rect 114058 278492 114074 278526
rect 111520 278480 114074 278492
rect 111520 278446 111536 278480
rect 112612 278446 112628 278480
rect 112744 278477 114074 278480
rect 112744 278460 114396 278477
rect 111452 278418 111486 278434
rect 111452 278274 111486 278290
rect 112662 278418 112696 278434
rect 112662 278274 112696 278290
rect 111520 278228 111536 278262
rect 112612 278228 112628 278262
rect 111334 278192 112628 278228
rect 111334 277868 111376 278192
rect 112744 278156 112780 278460
rect 113892 278441 114396 278460
rect 111520 278120 112780 278156
rect 112832 278382 113264 278416
rect 112832 278374 113012 278382
rect 112832 278120 112872 278374
rect 112996 278348 113012 278374
rect 114088 278348 114104 278382
rect 112928 278320 112962 278336
rect 112928 278256 112962 278272
rect 114138 278320 114172 278336
rect 114138 278256 114172 278272
rect 114324 278310 114396 278441
rect 112996 278216 113012 278244
rect 112994 278210 113012 278216
rect 114088 278216 114104 278244
rect 114324 278227 114342 278310
rect 114377 278227 114396 278310
rect 114088 278210 114274 278216
rect 112994 278170 114274 278210
rect 114324 278203 114396 278227
rect 111520 278086 111536 278120
rect 112612 278086 112628 278120
rect 112832 278084 113216 278120
rect 112832 278080 113012 278084
rect 111452 278058 111486 278074
rect 111452 277914 111486 277930
rect 112662 278058 112696 278074
rect 112832 278052 112872 278080
rect 112996 278050 113012 278080
rect 114088 278050 114104 278084
rect 112928 278022 112962 278038
rect 112928 277958 112962 277974
rect 114138 278022 114172 278038
rect 114138 277958 114172 277974
rect 112662 277914 112696 277930
rect 112996 277912 113012 277946
rect 114088 277912 114104 277946
rect 114234 277912 114274 278170
rect 111520 277868 111536 277902
rect 112612 277868 112628 277902
rect 111334 277832 112628 277868
rect 112994 277866 114455 277912
rect 113982 277759 114266 277764
rect 111312 277669 111328 277759
rect 114242 277669 114266 277759
rect 114652 279183 114862 279263
rect 114652 279149 114669 279183
rect 114845 279149 114862 279183
rect 114652 279148 114862 279149
rect 115027 279237 115178 279263
rect 114576 279121 114610 279137
rect 114576 278609 114610 278753
rect 114904 279121 114938 279137
rect 114653 278691 114669 278725
rect 114845 278691 114861 278725
rect 114904 278645 114938 278753
rect 114865 278628 114970 278645
rect 114865 278609 114885 278628
rect 114576 278561 114885 278609
rect 114576 278435 114610 278561
rect 114865 278560 114885 278561
rect 114948 278560 114970 278628
rect 114865 278538 114970 278560
rect 114653 278463 114669 278497
rect 114845 278463 114861 278497
rect 114576 278291 114610 278307
rect 114904 278435 114938 278538
rect 114904 278291 114938 278307
rect 114653 278245 114669 278279
rect 114845 278245 114861 278279
rect 114653 278208 114709 278245
rect 114805 278210 114861 278245
rect 114538 278169 114709 278208
rect 114804 278195 114991 278210
rect 114538 278043 114576 278169
rect 114804 278147 114868 278195
rect 114965 278147 114991 278195
rect 114804 278125 114991 278147
rect 114653 278055 114669 278089
rect 114845 278055 114861 278089
rect 114938 278043 114975 278125
rect 114538 278027 114610 278043
rect 114538 277899 114576 278027
rect 114538 277883 114610 277899
rect 114904 278027 114975 278043
rect 114938 277899 114975 278027
rect 114904 277883 114975 277899
rect 114653 277837 114669 277871
rect 114845 277837 114861 277871
rect 114455 277737 114489 277763
rect 114930 277763 115027 277821
rect 115061 277763 115144 279237
rect 115343 279183 115553 279263
rect 115343 279149 115360 279183
rect 115536 279149 115553 279183
rect 115343 279148 115553 279149
rect 115716 279237 115750 279263
rect 116183 279238 117169 279330
rect 115267 279121 115301 279137
rect 115267 278645 115301 278753
rect 115595 279121 115629 279137
rect 115344 278691 115360 278725
rect 115536 278691 115552 278725
rect 115235 278628 115340 278645
rect 115235 278560 115257 278628
rect 115320 278609 115340 278628
rect 115595 278609 115629 278753
rect 115320 278561 115629 278609
rect 115320 278560 115340 278561
rect 115235 278538 115340 278560
rect 115267 278435 115301 278538
rect 115344 278463 115360 278497
rect 115536 278463 115552 278497
rect 115267 278291 115301 278307
rect 115595 278435 115629 278561
rect 115595 278291 115629 278307
rect 115344 278245 115360 278279
rect 115536 278245 115552 278279
rect 115344 278210 115400 278245
rect 115214 278195 115401 278210
rect 115214 278147 115240 278195
rect 115337 278147 115401 278195
rect 115496 278208 115552 278245
rect 115496 278169 115667 278208
rect 115214 278125 115401 278147
rect 115230 278043 115267 278125
rect 115344 278055 115360 278089
rect 115536 278055 115552 278089
rect 115629 278043 115667 278169
rect 115230 278027 115301 278043
rect 115230 277899 115267 278027
rect 115230 277883 115301 277899
rect 115595 278027 115667 278043
rect 115629 277899 115667 278027
rect 115595 277883 115667 277899
rect 115344 277837 115360 277871
rect 115536 277837 115552 277871
rect 115178 277763 115275 277821
rect 114930 277737 115275 277763
rect 115959 279234 117169 279238
rect 115852 279233 117169 279234
rect 115852 279218 117239 279233
rect 115970 279208 117239 279218
rect 115970 279204 116147 279208
rect 115970 279100 115995 279204
rect 116131 279174 116147 279204
rect 117223 279174 117239 279208
rect 117391 279200 118685 279236
rect 115852 279084 115995 279100
rect 115959 278818 115995 279084
rect 116063 279146 116097 279162
rect 116063 278962 116097 278978
rect 117273 279146 117307 279162
rect 117273 278962 117307 278978
rect 116131 278916 116147 278950
rect 117223 278916 117239 278950
rect 117391 278916 117433 279200
rect 117577 279166 117593 279200
rect 118669 279166 118685 279200
rect 117509 279138 117543 279154
rect 117509 278994 117543 279010
rect 118719 279138 118753 279154
rect 118719 278994 118753 279010
rect 116131 278882 117433 278916
rect 117577 278948 117593 278982
rect 118669 278948 118685 278982
rect 117577 278912 118871 278948
rect 117373 278876 117433 278882
rect 117373 278840 118685 278876
rect 115959 278784 117239 278818
rect 116131 278750 116147 278784
rect 117223 278750 117239 278784
rect 116063 278722 116097 278738
rect 116063 278538 116097 278554
rect 117273 278722 117307 278738
rect 117273 278538 117307 278554
rect 116131 278492 116147 278526
rect 117223 278494 117239 278526
rect 117373 278516 117433 278840
rect 117577 278806 117593 278840
rect 118669 278806 118685 278840
rect 117509 278778 117543 278794
rect 117509 278634 117543 278650
rect 118719 278778 118753 278794
rect 118719 278634 118753 278650
rect 117577 278588 117593 278622
rect 118669 278588 118685 278622
rect 118829 278588 118871 278912
rect 117577 278552 118871 278588
rect 117373 278494 118685 278516
rect 117223 278492 118685 278494
rect 116131 278480 118685 278492
rect 116131 278477 117461 278480
rect 115809 278460 117461 278477
rect 115809 278441 116313 278460
rect 115809 278310 115881 278441
rect 116941 278382 117373 278416
rect 116101 278348 116117 278382
rect 117193 278374 117373 278382
rect 117193 278348 117209 278374
rect 115809 278227 115828 278310
rect 115863 278227 115881 278310
rect 116033 278320 116067 278336
rect 116033 278256 116067 278272
rect 117243 278320 117277 278336
rect 117243 278256 117277 278272
rect 115809 278203 115881 278227
rect 116101 278216 116117 278244
rect 115931 278210 116117 278216
rect 117193 278216 117209 278244
rect 117193 278210 117211 278216
rect 115931 278170 117211 278210
rect 115931 277912 115971 278170
rect 117333 278120 117373 278374
rect 117425 278156 117461 278460
rect 117577 278446 117593 278480
rect 118669 278446 118685 278480
rect 117509 278418 117543 278434
rect 117509 278274 117543 278290
rect 118719 278418 118753 278434
rect 118719 278274 118753 278290
rect 117577 278228 117593 278262
rect 118669 278228 118685 278262
rect 118829 278228 118871 278552
rect 117577 278192 118871 278228
rect 117425 278120 118685 278156
rect 116989 278084 117373 278120
rect 117577 278086 117593 278120
rect 118669 278086 118685 278120
rect 116101 278050 116117 278084
rect 117193 278080 117373 278084
rect 117193 278050 117209 278080
rect 117333 278052 117373 278080
rect 117509 278058 117543 278074
rect 116033 278022 116067 278038
rect 116033 277958 116067 277974
rect 117243 278022 117277 278038
rect 117243 277958 117277 277974
rect 116101 277912 116117 277946
rect 117193 277912 117209 277946
rect 117509 277914 117543 277930
rect 118719 278058 118753 278074
rect 118719 277914 118753 277930
rect 115750 277866 117211 277912
rect 117577 277868 117593 277902
rect 118669 277868 118685 277902
rect 118829 277868 118871 278192
rect 117577 277832 118871 277868
rect 115716 277737 115750 277763
rect 114455 277703 114515 277737
rect 115001 277703 115204 277737
rect 115690 277703 115750 277737
rect 115939 277759 116223 277764
rect 113036 277664 114266 277669
rect 113036 277572 114022 277664
rect 115061 277631 115144 277703
rect 115939 277669 115963 277759
rect 118877 277669 118893 277759
rect 115939 277664 117169 277669
rect 114455 277597 114515 277631
rect 115001 277597 115204 277631
rect 115690 277597 115750 277631
rect 111520 277534 112814 277570
rect 113036 277568 114246 277572
rect 114455 277571 114489 277597
rect 113036 277567 114353 277568
rect 111520 277500 111536 277534
rect 112612 277500 112628 277534
rect 111452 277472 111486 277488
rect 111452 277328 111486 277344
rect 112662 277472 112696 277488
rect 112662 277328 112696 277344
rect 111520 277282 111536 277316
rect 112612 277282 112628 277316
rect 111334 277246 112628 277282
rect 112772 277250 112814 277534
rect 112966 277552 114353 277567
rect 112966 277542 114235 277552
rect 112966 277508 112982 277542
rect 114058 277538 114235 277542
rect 114058 277508 114074 277538
rect 112898 277480 112932 277496
rect 112898 277296 112932 277312
rect 114108 277480 114142 277496
rect 114108 277296 114142 277312
rect 114210 277434 114235 277538
rect 114210 277418 114353 277434
rect 112966 277250 112982 277284
rect 114058 277250 114074 277284
rect 111334 276922 111376 277246
rect 112772 277216 114074 277250
rect 112772 277210 112832 277216
rect 111520 277174 112832 277210
rect 111520 277140 111536 277174
rect 112612 277140 112628 277174
rect 111452 277112 111486 277128
rect 111452 276968 111486 276984
rect 112662 277112 112696 277128
rect 112662 276968 112696 276984
rect 111520 276922 111536 276956
rect 112612 276922 112628 276956
rect 111334 276886 112628 276922
rect 111334 276562 111376 276886
rect 112772 276850 112832 277174
rect 114210 277152 114246 277418
rect 112966 277118 114246 277152
rect 112966 277084 112982 277118
rect 114058 277084 114074 277118
rect 112898 277056 112932 277072
rect 112898 276872 112932 276888
rect 114108 277056 114142 277072
rect 114108 276872 114142 276888
rect 111520 276828 112832 276850
rect 112966 276828 112982 276860
rect 111520 276826 112982 276828
rect 114058 276826 114074 276860
rect 111520 276814 114074 276826
rect 111520 276780 111536 276814
rect 112612 276780 112628 276814
rect 112744 276811 114074 276814
rect 112744 276794 114396 276811
rect 111452 276752 111486 276768
rect 111452 276608 111486 276624
rect 112662 276752 112696 276768
rect 112662 276608 112696 276624
rect 111520 276562 111536 276596
rect 112612 276562 112628 276596
rect 111334 276526 112628 276562
rect 111334 276202 111376 276526
rect 112744 276490 112780 276794
rect 113892 276775 114396 276794
rect 111520 276454 112780 276490
rect 112832 276716 113264 276750
rect 112832 276708 113012 276716
rect 112832 276454 112872 276708
rect 112996 276682 113012 276708
rect 114088 276682 114104 276716
rect 112928 276654 112962 276670
rect 112928 276590 112962 276606
rect 114138 276654 114172 276670
rect 114138 276590 114172 276606
rect 114324 276644 114396 276775
rect 112996 276550 113012 276578
rect 112994 276544 113012 276550
rect 114088 276550 114104 276578
rect 114324 276561 114342 276644
rect 114377 276561 114396 276644
rect 114088 276544 114274 276550
rect 112994 276504 114274 276544
rect 114324 276537 114396 276561
rect 111520 276420 111536 276454
rect 112612 276420 112628 276454
rect 112832 276418 113216 276454
rect 112832 276414 113012 276418
rect 111452 276392 111486 276408
rect 111452 276248 111486 276264
rect 112662 276392 112696 276408
rect 112832 276386 112872 276414
rect 112996 276384 113012 276414
rect 114088 276384 114104 276418
rect 112928 276356 112962 276372
rect 112928 276292 112962 276308
rect 114138 276356 114172 276372
rect 114138 276292 114172 276308
rect 112662 276248 112696 276264
rect 112996 276246 113012 276280
rect 114088 276246 114104 276280
rect 114234 276246 114274 276504
rect 111520 276202 111536 276236
rect 112612 276202 112628 276236
rect 111334 276166 112628 276202
rect 112994 276200 114455 276246
rect 113982 276093 114266 276098
rect 111312 276003 111328 276093
rect 114242 276003 114266 276093
rect 114652 277517 114862 277597
rect 114652 277483 114669 277517
rect 114845 277483 114862 277517
rect 114652 277482 114862 277483
rect 115027 277571 115178 277597
rect 114576 277455 114610 277471
rect 114576 276943 114610 277087
rect 114904 277455 114938 277471
rect 114653 277025 114669 277059
rect 114845 277025 114861 277059
rect 114904 276979 114938 277087
rect 114865 276962 114970 276979
rect 114865 276943 114885 276962
rect 114576 276895 114885 276943
rect 114576 276769 114610 276895
rect 114865 276894 114885 276895
rect 114948 276894 114970 276962
rect 114865 276872 114970 276894
rect 114653 276797 114669 276831
rect 114845 276797 114861 276831
rect 114576 276625 114610 276641
rect 114904 276769 114938 276872
rect 114904 276625 114938 276641
rect 114653 276579 114669 276613
rect 114845 276579 114861 276613
rect 114653 276542 114709 276579
rect 114805 276544 114861 276579
rect 114538 276503 114709 276542
rect 114804 276529 114991 276544
rect 114538 276377 114576 276503
rect 114804 276481 114868 276529
rect 114965 276481 114991 276529
rect 114804 276459 114991 276481
rect 114653 276389 114669 276423
rect 114845 276389 114861 276423
rect 114938 276377 114975 276459
rect 114538 276361 114610 276377
rect 114538 276233 114576 276361
rect 114538 276217 114610 276233
rect 114904 276361 114975 276377
rect 114938 276233 114975 276361
rect 114904 276217 114975 276233
rect 114653 276171 114669 276205
rect 114845 276171 114861 276205
rect 114455 276071 114489 276097
rect 114930 276097 115027 276155
rect 115061 276097 115144 277571
rect 115343 277517 115553 277597
rect 115343 277483 115360 277517
rect 115536 277483 115553 277517
rect 115343 277482 115553 277483
rect 115716 277571 115750 277597
rect 116183 277572 117169 277664
rect 115267 277455 115301 277471
rect 115267 276979 115301 277087
rect 115595 277455 115629 277471
rect 115344 277025 115360 277059
rect 115536 277025 115552 277059
rect 115235 276962 115340 276979
rect 115235 276894 115257 276962
rect 115320 276943 115340 276962
rect 115595 276943 115629 277087
rect 115320 276895 115629 276943
rect 115320 276894 115340 276895
rect 115235 276872 115340 276894
rect 115267 276769 115301 276872
rect 115344 276797 115360 276831
rect 115536 276797 115552 276831
rect 115267 276625 115301 276641
rect 115595 276769 115629 276895
rect 115595 276625 115629 276641
rect 115344 276579 115360 276613
rect 115536 276579 115552 276613
rect 115344 276544 115400 276579
rect 115214 276529 115401 276544
rect 115214 276481 115240 276529
rect 115337 276481 115401 276529
rect 115496 276542 115552 276579
rect 115496 276503 115667 276542
rect 115214 276459 115401 276481
rect 115230 276377 115267 276459
rect 115344 276389 115360 276423
rect 115536 276389 115552 276423
rect 115629 276377 115667 276503
rect 115230 276361 115301 276377
rect 115230 276233 115267 276361
rect 115230 276217 115301 276233
rect 115595 276361 115667 276377
rect 115629 276233 115667 276361
rect 115595 276217 115667 276233
rect 115344 276171 115360 276205
rect 115536 276171 115552 276205
rect 115178 276097 115275 276155
rect 114930 276071 115275 276097
rect 115959 277568 117169 277572
rect 115852 277567 117169 277568
rect 115852 277552 117239 277567
rect 115970 277542 117239 277552
rect 115970 277538 116147 277542
rect 115970 277434 115995 277538
rect 116131 277508 116147 277538
rect 117223 277508 117239 277542
rect 117391 277534 118685 277570
rect 115852 277418 115995 277434
rect 115959 277152 115995 277418
rect 116063 277480 116097 277496
rect 116063 277296 116097 277312
rect 117273 277480 117307 277496
rect 117273 277296 117307 277312
rect 116131 277250 116147 277284
rect 117223 277250 117239 277284
rect 117391 277250 117433 277534
rect 117577 277500 117593 277534
rect 118669 277500 118685 277534
rect 117509 277472 117543 277488
rect 117509 277328 117543 277344
rect 118719 277472 118753 277488
rect 118719 277328 118753 277344
rect 116131 277216 117433 277250
rect 117577 277282 117593 277316
rect 118669 277282 118685 277316
rect 117577 277246 118871 277282
rect 117373 277210 117433 277216
rect 117373 277174 118685 277210
rect 115959 277118 117239 277152
rect 116131 277084 116147 277118
rect 117223 277084 117239 277118
rect 116063 277056 116097 277072
rect 116063 276872 116097 276888
rect 117273 277056 117307 277072
rect 117273 276872 117307 276888
rect 116131 276826 116147 276860
rect 117223 276828 117239 276860
rect 117373 276850 117433 277174
rect 117577 277140 117593 277174
rect 118669 277140 118685 277174
rect 117509 277112 117543 277128
rect 117509 276968 117543 276984
rect 118719 277112 118753 277128
rect 118719 276968 118753 276984
rect 117577 276922 117593 276956
rect 118669 276922 118685 276956
rect 118829 276922 118871 277246
rect 117577 276886 118871 276922
rect 117373 276828 118685 276850
rect 117223 276826 118685 276828
rect 116131 276814 118685 276826
rect 116131 276811 117461 276814
rect 115809 276794 117461 276811
rect 115809 276775 116313 276794
rect 115809 276644 115881 276775
rect 116941 276716 117373 276750
rect 116101 276682 116117 276716
rect 117193 276708 117373 276716
rect 117193 276682 117209 276708
rect 115809 276561 115828 276644
rect 115863 276561 115881 276644
rect 116033 276654 116067 276670
rect 116033 276590 116067 276606
rect 117243 276654 117277 276670
rect 117243 276590 117277 276606
rect 115809 276537 115881 276561
rect 116101 276550 116117 276578
rect 115931 276544 116117 276550
rect 117193 276550 117209 276578
rect 117193 276544 117211 276550
rect 115931 276504 117211 276544
rect 115931 276246 115971 276504
rect 117333 276454 117373 276708
rect 117425 276490 117461 276794
rect 117577 276780 117593 276814
rect 118669 276780 118685 276814
rect 117509 276752 117543 276768
rect 117509 276608 117543 276624
rect 118719 276752 118753 276768
rect 118719 276608 118753 276624
rect 117577 276562 117593 276596
rect 118669 276562 118685 276596
rect 118829 276562 118871 276886
rect 117577 276526 118871 276562
rect 117425 276454 118685 276490
rect 116989 276418 117373 276454
rect 117577 276420 117593 276454
rect 118669 276420 118685 276454
rect 116101 276384 116117 276418
rect 117193 276414 117373 276418
rect 117193 276384 117209 276414
rect 117333 276386 117373 276414
rect 117509 276392 117543 276408
rect 116033 276356 116067 276372
rect 116033 276292 116067 276308
rect 117243 276356 117277 276372
rect 117243 276292 117277 276308
rect 116101 276246 116117 276280
rect 117193 276246 117209 276280
rect 117509 276248 117543 276264
rect 118719 276392 118753 276408
rect 118719 276248 118753 276264
rect 115750 276200 117211 276246
rect 117577 276202 117593 276236
rect 118669 276202 118685 276236
rect 118829 276202 118871 276526
rect 117577 276166 118871 276202
rect 115716 276071 115750 276097
rect 114455 276037 114515 276071
rect 115001 276037 115204 276071
rect 115690 276037 115750 276071
rect 115939 276093 116223 276098
rect 113036 275998 114266 276003
rect 113036 275906 114022 275998
rect 115061 275965 115144 276037
rect 115939 276003 115963 276093
rect 118877 276003 118893 276093
rect 115939 275998 117169 276003
rect 114455 275931 114515 275965
rect 115001 275931 115204 275965
rect 115690 275931 115750 275965
rect 111520 275868 112814 275904
rect 113036 275902 114246 275906
rect 114455 275905 114489 275931
rect 113036 275901 114353 275902
rect 111520 275834 111536 275868
rect 112612 275834 112628 275868
rect 111452 275806 111486 275822
rect 111452 275662 111486 275678
rect 112662 275806 112696 275822
rect 112662 275662 112696 275678
rect 111520 275616 111536 275650
rect 112612 275616 112628 275650
rect 111334 275580 112628 275616
rect 112772 275584 112814 275868
rect 112966 275886 114353 275901
rect 112966 275876 114235 275886
rect 112966 275842 112982 275876
rect 114058 275872 114235 275876
rect 114058 275842 114074 275872
rect 112898 275814 112932 275830
rect 112898 275630 112932 275646
rect 114108 275814 114142 275830
rect 114108 275630 114142 275646
rect 114210 275768 114235 275872
rect 114210 275752 114353 275768
rect 112966 275584 112982 275618
rect 114058 275584 114074 275618
rect 111334 275256 111376 275580
rect 112772 275550 114074 275584
rect 112772 275544 112832 275550
rect 111520 275508 112832 275544
rect 111520 275474 111536 275508
rect 112612 275474 112628 275508
rect 111452 275446 111486 275462
rect 111452 275302 111486 275318
rect 112662 275446 112696 275462
rect 112662 275302 112696 275318
rect 111520 275256 111536 275290
rect 112612 275256 112628 275290
rect 111334 275220 112628 275256
rect 111334 274896 111376 275220
rect 112772 275184 112832 275508
rect 114210 275486 114246 275752
rect 112966 275452 114246 275486
rect 112966 275418 112982 275452
rect 114058 275418 114074 275452
rect 112898 275390 112932 275406
rect 112898 275206 112932 275222
rect 114108 275390 114142 275406
rect 114108 275206 114142 275222
rect 111520 275162 112832 275184
rect 112966 275162 112982 275194
rect 111520 275160 112982 275162
rect 114058 275160 114074 275194
rect 111520 275148 114074 275160
rect 111520 275114 111536 275148
rect 112612 275114 112628 275148
rect 112744 275145 114074 275148
rect 112744 275128 114396 275145
rect 111452 275086 111486 275102
rect 111452 274942 111486 274958
rect 112662 275086 112696 275102
rect 112662 274942 112696 274958
rect 111520 274896 111536 274930
rect 112612 274896 112628 274930
rect 111334 274860 112628 274896
rect 111334 274536 111376 274860
rect 112744 274824 112780 275128
rect 113892 275109 114396 275128
rect 111520 274788 112780 274824
rect 112832 275050 113264 275084
rect 112832 275042 113012 275050
rect 112832 274788 112872 275042
rect 112996 275016 113012 275042
rect 114088 275016 114104 275050
rect 112928 274988 112962 275004
rect 112928 274924 112962 274940
rect 114138 274988 114172 275004
rect 114138 274924 114172 274940
rect 114324 274978 114396 275109
rect 112996 274884 113012 274912
rect 112994 274878 113012 274884
rect 114088 274884 114104 274912
rect 114324 274895 114342 274978
rect 114377 274895 114396 274978
rect 114088 274878 114274 274884
rect 112994 274838 114274 274878
rect 114324 274871 114396 274895
rect 111520 274754 111536 274788
rect 112612 274754 112628 274788
rect 112832 274752 113216 274788
rect 112832 274748 113012 274752
rect 111452 274726 111486 274742
rect 111452 274582 111486 274598
rect 112662 274726 112696 274742
rect 112832 274720 112872 274748
rect 112996 274718 113012 274748
rect 114088 274718 114104 274752
rect 112928 274690 112962 274706
rect 112928 274626 112962 274642
rect 114138 274690 114172 274706
rect 114138 274626 114172 274642
rect 112662 274582 112696 274598
rect 112996 274580 113012 274614
rect 114088 274580 114104 274614
rect 114234 274580 114274 274838
rect 111520 274536 111536 274570
rect 112612 274536 112628 274570
rect 111334 274500 112628 274536
rect 112994 274534 114455 274580
rect 113982 274427 114266 274432
rect 111312 274337 111328 274427
rect 114242 274337 114266 274427
rect 114652 275851 114862 275931
rect 114652 275817 114669 275851
rect 114845 275817 114862 275851
rect 114652 275816 114862 275817
rect 115027 275905 115178 275931
rect 114576 275789 114610 275805
rect 114576 275277 114610 275421
rect 114904 275789 114938 275805
rect 114653 275359 114669 275393
rect 114845 275359 114861 275393
rect 114904 275313 114938 275421
rect 114865 275296 114970 275313
rect 114865 275277 114885 275296
rect 114576 275229 114885 275277
rect 114576 275103 114610 275229
rect 114865 275228 114885 275229
rect 114948 275228 114970 275296
rect 114865 275206 114970 275228
rect 114653 275131 114669 275165
rect 114845 275131 114861 275165
rect 114576 274959 114610 274975
rect 114904 275103 114938 275206
rect 114904 274959 114938 274975
rect 114653 274913 114669 274947
rect 114845 274913 114861 274947
rect 114653 274876 114709 274913
rect 114805 274878 114861 274913
rect 114538 274837 114709 274876
rect 114804 274863 114991 274878
rect 114538 274711 114576 274837
rect 114804 274815 114868 274863
rect 114965 274815 114991 274863
rect 114804 274793 114991 274815
rect 114653 274723 114669 274757
rect 114845 274723 114861 274757
rect 114938 274711 114975 274793
rect 114538 274695 114610 274711
rect 114538 274567 114576 274695
rect 114538 274551 114610 274567
rect 114904 274695 114975 274711
rect 114938 274567 114975 274695
rect 114904 274551 114975 274567
rect 114653 274505 114669 274539
rect 114845 274505 114861 274539
rect 114455 274405 114489 274431
rect 114930 274431 115027 274489
rect 115061 274431 115144 275905
rect 115343 275851 115553 275931
rect 115343 275817 115360 275851
rect 115536 275817 115553 275851
rect 115343 275816 115553 275817
rect 115716 275905 115750 275931
rect 116183 275906 117169 275998
rect 115267 275789 115301 275805
rect 115267 275313 115301 275421
rect 115595 275789 115629 275805
rect 115344 275359 115360 275393
rect 115536 275359 115552 275393
rect 115235 275296 115340 275313
rect 115235 275228 115257 275296
rect 115320 275277 115340 275296
rect 115595 275277 115629 275421
rect 115320 275229 115629 275277
rect 115320 275228 115340 275229
rect 115235 275206 115340 275228
rect 115267 275103 115301 275206
rect 115344 275131 115360 275165
rect 115536 275131 115552 275165
rect 115267 274959 115301 274975
rect 115595 275103 115629 275229
rect 115595 274959 115629 274975
rect 115344 274913 115360 274947
rect 115536 274913 115552 274947
rect 115344 274878 115400 274913
rect 115214 274863 115401 274878
rect 115214 274815 115240 274863
rect 115337 274815 115401 274863
rect 115496 274876 115552 274913
rect 115496 274837 115667 274876
rect 115214 274793 115401 274815
rect 115230 274711 115267 274793
rect 115344 274723 115360 274757
rect 115536 274723 115552 274757
rect 115629 274711 115667 274837
rect 115230 274695 115301 274711
rect 115230 274567 115267 274695
rect 115230 274551 115301 274567
rect 115595 274695 115667 274711
rect 115629 274567 115667 274695
rect 115595 274551 115667 274567
rect 115344 274505 115360 274539
rect 115536 274505 115552 274539
rect 115178 274431 115275 274489
rect 114930 274405 115275 274431
rect 115959 275902 117169 275906
rect 115852 275901 117169 275902
rect 115852 275886 117239 275901
rect 115970 275876 117239 275886
rect 115970 275872 116147 275876
rect 115970 275768 115995 275872
rect 116131 275842 116147 275872
rect 117223 275842 117239 275876
rect 117391 275868 118685 275904
rect 115852 275752 115995 275768
rect 115959 275486 115995 275752
rect 116063 275814 116097 275830
rect 116063 275630 116097 275646
rect 117273 275814 117307 275830
rect 117273 275630 117307 275646
rect 116131 275584 116147 275618
rect 117223 275584 117239 275618
rect 117391 275584 117433 275868
rect 117577 275834 117593 275868
rect 118669 275834 118685 275868
rect 117509 275806 117543 275822
rect 117509 275662 117543 275678
rect 118719 275806 118753 275822
rect 118719 275662 118753 275678
rect 116131 275550 117433 275584
rect 117577 275616 117593 275650
rect 118669 275616 118685 275650
rect 117577 275580 118871 275616
rect 117373 275544 117433 275550
rect 117373 275508 118685 275544
rect 115959 275452 117239 275486
rect 116131 275418 116147 275452
rect 117223 275418 117239 275452
rect 116063 275390 116097 275406
rect 116063 275206 116097 275222
rect 117273 275390 117307 275406
rect 117273 275206 117307 275222
rect 116131 275160 116147 275194
rect 117223 275162 117239 275194
rect 117373 275184 117433 275508
rect 117577 275474 117593 275508
rect 118669 275474 118685 275508
rect 117509 275446 117543 275462
rect 117509 275302 117543 275318
rect 118719 275446 118753 275462
rect 118719 275302 118753 275318
rect 117577 275256 117593 275290
rect 118669 275256 118685 275290
rect 118829 275256 118871 275580
rect 117577 275220 118871 275256
rect 117373 275162 118685 275184
rect 117223 275160 118685 275162
rect 116131 275148 118685 275160
rect 116131 275145 117461 275148
rect 115809 275128 117461 275145
rect 115809 275109 116313 275128
rect 115809 274978 115881 275109
rect 116941 275050 117373 275084
rect 116101 275016 116117 275050
rect 117193 275042 117373 275050
rect 117193 275016 117209 275042
rect 115809 274895 115828 274978
rect 115863 274895 115881 274978
rect 116033 274988 116067 275004
rect 116033 274924 116067 274940
rect 117243 274988 117277 275004
rect 117243 274924 117277 274940
rect 115809 274871 115881 274895
rect 116101 274884 116117 274912
rect 115931 274878 116117 274884
rect 117193 274884 117209 274912
rect 117193 274878 117211 274884
rect 115931 274838 117211 274878
rect 115931 274580 115971 274838
rect 117333 274788 117373 275042
rect 117425 274824 117461 275128
rect 117577 275114 117593 275148
rect 118669 275114 118685 275148
rect 117509 275086 117543 275102
rect 117509 274942 117543 274958
rect 118719 275086 118753 275102
rect 118719 274942 118753 274958
rect 117577 274896 117593 274930
rect 118669 274896 118685 274930
rect 118829 274896 118871 275220
rect 117577 274860 118871 274896
rect 117425 274788 118685 274824
rect 116989 274752 117373 274788
rect 117577 274754 117593 274788
rect 118669 274754 118685 274788
rect 116101 274718 116117 274752
rect 117193 274748 117373 274752
rect 117193 274718 117209 274748
rect 117333 274720 117373 274748
rect 117509 274726 117543 274742
rect 116033 274690 116067 274706
rect 116033 274626 116067 274642
rect 117243 274690 117277 274706
rect 117243 274626 117277 274642
rect 116101 274580 116117 274614
rect 117193 274580 117209 274614
rect 117509 274582 117543 274598
rect 118719 274726 118753 274742
rect 118719 274582 118753 274598
rect 115750 274534 117211 274580
rect 117577 274536 117593 274570
rect 118669 274536 118685 274570
rect 118829 274536 118871 274860
rect 117577 274500 118871 274536
rect 115716 274405 115750 274431
rect 114455 274371 114515 274405
rect 115001 274371 115204 274405
rect 115690 274371 115750 274405
rect 115939 274427 116223 274432
rect 113036 274332 114266 274337
rect 113036 274240 114022 274332
rect 115061 274299 115144 274371
rect 115939 274337 115963 274427
rect 118877 274337 118893 274427
rect 115939 274332 117169 274337
rect 114455 274265 114515 274299
rect 115001 274265 115204 274299
rect 115690 274265 115750 274299
rect 111520 274202 112814 274238
rect 113036 274236 114246 274240
rect 114455 274239 114489 274265
rect 113036 274235 114353 274236
rect 111520 274168 111536 274202
rect 112612 274168 112628 274202
rect 111452 274140 111486 274156
rect 111452 273996 111486 274012
rect 112662 274140 112696 274156
rect 112662 273996 112696 274012
rect 111520 273950 111536 273984
rect 112612 273950 112628 273984
rect 111334 273914 112628 273950
rect 112772 273918 112814 274202
rect 112966 274220 114353 274235
rect 112966 274210 114235 274220
rect 112966 274176 112982 274210
rect 114058 274206 114235 274210
rect 114058 274176 114074 274206
rect 112898 274148 112932 274164
rect 112898 273964 112932 273980
rect 114108 274148 114142 274164
rect 114108 273964 114142 273980
rect 114210 274102 114235 274206
rect 114210 274086 114353 274102
rect 112966 273918 112982 273952
rect 114058 273918 114074 273952
rect 111334 273590 111376 273914
rect 112772 273884 114074 273918
rect 112772 273878 112832 273884
rect 111520 273842 112832 273878
rect 111520 273808 111536 273842
rect 112612 273808 112628 273842
rect 111452 273780 111486 273796
rect 111452 273636 111486 273652
rect 112662 273780 112696 273796
rect 112662 273636 112696 273652
rect 111520 273590 111536 273624
rect 112612 273590 112628 273624
rect 111334 273554 112628 273590
rect 111334 273230 111376 273554
rect 112772 273518 112832 273842
rect 114210 273820 114246 274086
rect 112966 273786 114246 273820
rect 112966 273752 112982 273786
rect 114058 273752 114074 273786
rect 112898 273724 112932 273740
rect 112898 273540 112932 273556
rect 114108 273724 114142 273740
rect 114108 273540 114142 273556
rect 111520 273496 112832 273518
rect 112966 273496 112982 273528
rect 111520 273494 112982 273496
rect 114058 273494 114074 273528
rect 111520 273482 114074 273494
rect 111520 273448 111536 273482
rect 112612 273448 112628 273482
rect 112744 273479 114074 273482
rect 112744 273462 114396 273479
rect 111452 273420 111486 273436
rect 111452 273276 111486 273292
rect 112662 273420 112696 273436
rect 112662 273276 112696 273292
rect 111520 273230 111536 273264
rect 112612 273230 112628 273264
rect 111334 273194 112628 273230
rect 111334 272870 111376 273194
rect 112744 273158 112780 273462
rect 113892 273443 114396 273462
rect 111520 273122 112780 273158
rect 112832 273384 113264 273418
rect 112832 273376 113012 273384
rect 112832 273122 112872 273376
rect 112996 273350 113012 273376
rect 114088 273350 114104 273384
rect 112928 273322 112962 273338
rect 112928 273258 112962 273274
rect 114138 273322 114172 273338
rect 114138 273258 114172 273274
rect 114324 273312 114396 273443
rect 112996 273218 113012 273246
rect 112994 273212 113012 273218
rect 114088 273218 114104 273246
rect 114324 273229 114342 273312
rect 114377 273229 114396 273312
rect 114088 273212 114274 273218
rect 112994 273172 114274 273212
rect 114324 273205 114396 273229
rect 111520 273088 111536 273122
rect 112612 273088 112628 273122
rect 112832 273086 113216 273122
rect 112832 273082 113012 273086
rect 111452 273060 111486 273076
rect 111452 272916 111486 272932
rect 112662 273060 112696 273076
rect 112832 273054 112872 273082
rect 112996 273052 113012 273082
rect 114088 273052 114104 273086
rect 112928 273024 112962 273040
rect 112928 272960 112962 272976
rect 114138 273024 114172 273040
rect 114138 272960 114172 272976
rect 112662 272916 112696 272932
rect 112996 272914 113012 272948
rect 114088 272914 114104 272948
rect 114234 272914 114274 273172
rect 111520 272870 111536 272904
rect 112612 272870 112628 272904
rect 111334 272834 112628 272870
rect 112994 272868 114455 272914
rect 113982 272761 114266 272766
rect 111046 272683 111200 272699
rect 111312 272671 111328 272761
rect 114242 272671 114266 272761
rect 114652 274185 114862 274265
rect 114652 274151 114669 274185
rect 114845 274151 114862 274185
rect 114652 274150 114862 274151
rect 115027 274239 115178 274265
rect 114576 274123 114610 274139
rect 114576 273611 114610 273755
rect 114904 274123 114938 274139
rect 114653 273693 114669 273727
rect 114845 273693 114861 273727
rect 114904 273647 114938 273755
rect 114865 273630 114970 273647
rect 114865 273611 114885 273630
rect 114576 273563 114885 273611
rect 114576 273437 114610 273563
rect 114865 273562 114885 273563
rect 114948 273562 114970 273630
rect 114865 273540 114970 273562
rect 114653 273465 114669 273499
rect 114845 273465 114861 273499
rect 114576 273293 114610 273309
rect 114904 273437 114938 273540
rect 114904 273293 114938 273309
rect 114653 273247 114669 273281
rect 114845 273247 114861 273281
rect 114653 273210 114709 273247
rect 114805 273212 114861 273247
rect 114538 273171 114709 273210
rect 114804 273197 114991 273212
rect 114538 273045 114576 273171
rect 114804 273149 114868 273197
rect 114965 273149 114991 273197
rect 114804 273127 114991 273149
rect 114653 273057 114669 273091
rect 114845 273057 114861 273091
rect 114938 273045 114975 273127
rect 114538 273029 114610 273045
rect 114538 272901 114576 273029
rect 114538 272885 114610 272901
rect 114904 273029 114975 273045
rect 114938 272901 114975 273029
rect 114904 272885 114975 272901
rect 114653 272839 114669 272873
rect 114845 272839 114861 272873
rect 114455 272739 114489 272765
rect 114928 272793 115027 272825
rect 115061 272793 115144 274239
rect 115343 274185 115553 274265
rect 115343 274151 115360 274185
rect 115536 274151 115553 274185
rect 115343 274150 115553 274151
rect 115716 274239 115750 274265
rect 116183 274240 117169 274332
rect 115267 274123 115301 274139
rect 115267 273647 115301 273755
rect 115595 274123 115629 274139
rect 115344 273693 115360 273727
rect 115536 273693 115552 273727
rect 115235 273630 115340 273647
rect 115235 273562 115257 273630
rect 115320 273611 115340 273630
rect 115595 273611 115629 273755
rect 115320 273563 115629 273611
rect 115320 273562 115340 273563
rect 115235 273540 115340 273562
rect 115267 273437 115301 273540
rect 115344 273465 115360 273499
rect 115536 273465 115552 273499
rect 115267 273293 115301 273309
rect 115595 273437 115629 273563
rect 115595 273293 115629 273309
rect 115344 273247 115360 273281
rect 115536 273247 115552 273281
rect 115344 273212 115400 273247
rect 115214 273197 115401 273212
rect 115214 273149 115240 273197
rect 115337 273149 115401 273197
rect 115496 273210 115552 273247
rect 115496 273171 115667 273210
rect 115214 273127 115401 273149
rect 115230 273045 115267 273127
rect 115344 273057 115360 273091
rect 115536 273057 115552 273091
rect 115629 273045 115667 273171
rect 115230 273029 115301 273045
rect 115230 272901 115267 273029
rect 115230 272885 115301 272901
rect 115595 273029 115667 273045
rect 115629 272901 115667 273029
rect 115595 272885 115667 272901
rect 115344 272839 115360 272873
rect 115536 272839 115552 272873
rect 115178 272793 115275 272825
rect 114928 272739 114982 272793
rect 115228 272739 115275 272793
rect 115959 274236 117169 274240
rect 115852 274235 117169 274236
rect 115852 274220 117239 274235
rect 115970 274210 117239 274220
rect 115970 274206 116147 274210
rect 115970 274102 115995 274206
rect 116131 274176 116147 274206
rect 117223 274176 117239 274210
rect 117391 274202 118685 274238
rect 115852 274086 115995 274102
rect 115959 273820 115995 274086
rect 116063 274148 116097 274164
rect 116063 273964 116097 273980
rect 117273 274148 117307 274164
rect 117273 273964 117307 273980
rect 116131 273918 116147 273952
rect 117223 273918 117239 273952
rect 117391 273918 117433 274202
rect 117577 274168 117593 274202
rect 118669 274168 118685 274202
rect 117509 274140 117543 274156
rect 117509 273996 117543 274012
rect 118719 274140 118753 274156
rect 118719 273996 118753 274012
rect 116131 273884 117433 273918
rect 117577 273950 117593 273984
rect 118669 273950 118685 273984
rect 117577 273914 118871 273950
rect 117373 273878 117433 273884
rect 117373 273842 118685 273878
rect 115959 273786 117239 273820
rect 116131 273752 116147 273786
rect 117223 273752 117239 273786
rect 116063 273724 116097 273740
rect 116063 273540 116097 273556
rect 117273 273724 117307 273740
rect 117273 273540 117307 273556
rect 116131 273494 116147 273528
rect 117223 273496 117239 273528
rect 117373 273518 117433 273842
rect 117577 273808 117593 273842
rect 118669 273808 118685 273842
rect 117509 273780 117543 273796
rect 117509 273636 117543 273652
rect 118719 273780 118753 273796
rect 118719 273636 118753 273652
rect 117577 273590 117593 273624
rect 118669 273590 118685 273624
rect 118829 273590 118871 273914
rect 117577 273554 118871 273590
rect 117373 273496 118685 273518
rect 117223 273494 118685 273496
rect 116131 273482 118685 273494
rect 116131 273479 117461 273482
rect 115809 273462 117461 273479
rect 115809 273443 116313 273462
rect 115809 273312 115881 273443
rect 116941 273384 117373 273418
rect 116101 273350 116117 273384
rect 117193 273376 117373 273384
rect 117193 273350 117209 273376
rect 115809 273229 115828 273312
rect 115863 273229 115881 273312
rect 116033 273322 116067 273338
rect 116033 273258 116067 273274
rect 117243 273322 117277 273338
rect 117243 273258 117277 273274
rect 115809 273205 115881 273229
rect 116101 273218 116117 273246
rect 115931 273212 116117 273218
rect 117193 273218 117209 273246
rect 117193 273212 117211 273218
rect 115931 273172 117211 273212
rect 115931 272914 115971 273172
rect 117333 273122 117373 273376
rect 117425 273158 117461 273462
rect 117577 273448 117593 273482
rect 118669 273448 118685 273482
rect 117509 273420 117543 273436
rect 117509 273276 117543 273292
rect 118719 273420 118753 273436
rect 118719 273276 118753 273292
rect 117577 273230 117593 273264
rect 118669 273230 118685 273264
rect 118829 273230 118871 273554
rect 117577 273194 118871 273230
rect 117425 273122 118685 273158
rect 116989 273086 117373 273122
rect 117577 273088 117593 273122
rect 118669 273088 118685 273122
rect 116101 273052 116117 273086
rect 117193 273082 117373 273086
rect 117193 273052 117209 273082
rect 117333 273054 117373 273082
rect 117509 273060 117543 273076
rect 116033 273024 116067 273040
rect 116033 272960 116067 272976
rect 117243 273024 117277 273040
rect 117243 272960 117277 272976
rect 116101 272914 116117 272948
rect 117193 272914 117209 272948
rect 117509 272916 117543 272932
rect 118719 273060 118753 273076
rect 118719 272916 118753 272932
rect 115750 272868 117211 272914
rect 117577 272870 117593 272904
rect 118669 272870 118685 272904
rect 118829 272870 118871 273194
rect 117577 272834 118871 272870
rect 115716 272739 115750 272765
rect 114455 272705 114515 272739
rect 115690 272705 115750 272739
rect 115939 272761 116223 272766
rect 118762 272761 119005 272762
rect 109967 270177 110259 270193
rect 106281 270169 110259 270177
rect 111939 272249 112069 272265
rect 112673 272249 113101 272671
rect 113982 272666 114266 272671
rect 114928 272417 114982 272705
rect 115228 272417 115275 272705
rect 115939 272671 115963 272761
rect 118877 272699 119005 272761
rect 118877 272683 119159 272699
rect 119938 281067 120227 281165
rect 118877 272671 119158 272683
rect 115939 272666 116223 272671
rect 114928 272372 115275 272417
rect 116523 272249 119158 272671
rect 107329 268607 108364 270169
rect 112069 272125 112167 272249
rect 118956 272125 119021 272249
rect 116590 272098 118192 272125
rect 113800 272014 114102 272051
rect 113800 271699 113840 272014
rect 114065 271699 114102 272014
rect 114984 272036 115601 272048
rect 114984 272016 118841 272036
rect 114984 271918 115017 272016
rect 115559 271996 118841 272016
rect 115559 271981 115897 271996
rect 115559 271918 115601 271981
rect 114984 271886 115601 271918
rect 113800 271668 114102 271699
rect 112307 271634 112367 271668
rect 114150 271634 114210 271668
rect 112307 271608 112341 271634
rect 113068 271629 113461 271634
rect 113068 271540 113091 271629
rect 113431 271540 113461 271629
rect 113068 271524 113461 271540
rect 114176 271608 114210 271634
rect 112578 271353 112594 271387
rect 112722 271353 112994 271387
rect 113122 271353 113394 271387
rect 113522 271353 113794 271387
rect 113922 271353 113938 271387
rect 112532 271294 112566 271310
rect 112532 271102 112566 271118
rect 112750 271294 112784 271310
rect 112750 271102 112784 271118
rect 112838 271059 112886 271353
rect 112932 271294 112966 271310
rect 112932 271102 112966 271118
rect 113150 271294 113184 271310
rect 113150 271102 113184 271118
rect 113332 271294 113366 271310
rect 113332 271102 113366 271118
rect 113550 271294 113584 271310
rect 113550 271102 113584 271118
rect 113634 271059 113682 271353
rect 113732 271294 113766 271310
rect 113732 271102 113766 271118
rect 113950 271294 113984 271310
rect 113950 271102 113984 271118
rect 112578 271025 112594 271059
rect 112722 271025 112994 271059
rect 113122 271025 113394 271059
rect 113522 271025 113794 271059
rect 113922 271025 113938 271059
rect 112307 270817 112341 270843
rect 114329 271567 114389 271588
rect 114210 271554 114389 271567
rect 115443 271554 115503 271588
rect 114210 271528 114363 271554
rect 114210 270843 114329 271528
rect 114176 270832 114329 270843
rect 114637 271324 114653 271358
rect 114781 271324 114797 271358
rect 114591 271265 114625 271281
rect 114591 271073 114625 271089
rect 114809 271279 114843 271281
rect 114890 271279 114942 271554
rect 115469 271528 115503 271554
rect 115337 271373 115382 271375
rect 115060 271358 115382 271373
rect 115037 271324 115053 271358
rect 115181 271331 115382 271358
rect 115181 271324 115197 271331
rect 114991 271279 115025 271281
rect 114809 271265 115025 271279
rect 114843 271229 114991 271265
rect 114809 271073 114843 271089
rect 114991 271073 115025 271089
rect 115209 271265 115243 271281
rect 115209 271073 115243 271089
rect 114637 270996 114653 271030
rect 114781 270996 115053 271030
rect 115181 271014 115197 271030
rect 115337 271014 115382 271331
rect 115181 270996 115382 271014
rect 115074 270973 115382 270996
rect 115074 270972 115369 270973
rect 114176 270817 114363 270832
rect 112307 270783 112367 270817
rect 114150 270806 114363 270817
rect 115469 270806 115503 270832
rect 114150 270789 114389 270806
rect 114150 270783 114210 270789
rect 114329 270772 114389 270789
rect 115443 270772 115503 270806
rect 115648 270763 115700 271981
rect 115881 271962 115897 271981
rect 116025 271962 116297 271996
rect 116425 271962 116697 271996
rect 116825 271962 117097 271996
rect 117225 271962 117497 271996
rect 117625 271962 117897 271996
rect 118025 271962 118297 271996
rect 118425 271962 118697 271996
rect 118825 271962 118841 271996
rect 115835 271912 115869 271928
rect 115835 270820 115869 270836
rect 116053 271912 116087 271928
rect 116053 270820 116087 270836
rect 116235 271912 116269 271928
rect 116235 270820 116269 270836
rect 116453 271912 116487 271928
rect 116453 270820 116487 270836
rect 116635 271912 116669 271928
rect 116635 270820 116669 270836
rect 116853 271912 116887 271928
rect 116853 270820 116887 270836
rect 117035 271912 117069 271928
rect 117035 270820 117069 270836
rect 117253 271912 117287 271928
rect 117253 270820 117287 270836
rect 117435 271912 117469 271928
rect 117435 270820 117469 270836
rect 117653 271912 117687 271928
rect 117653 270820 117687 270836
rect 117835 271912 117869 271928
rect 117835 270820 117869 270836
rect 118053 271912 118087 271928
rect 118053 270820 118087 270836
rect 118235 271912 118269 271928
rect 118235 270820 118269 270836
rect 118453 271912 118487 271928
rect 118453 270820 118487 270836
rect 118635 271912 118669 271928
rect 118635 270820 118669 270836
rect 118853 271912 118887 271928
rect 118853 270820 118887 270836
rect 115881 270763 115897 270786
rect 115648 270752 115897 270763
rect 116025 270752 116297 270786
rect 116425 270752 116697 270786
rect 116825 270752 117097 270786
rect 117225 270752 117497 270786
rect 117625 270752 117897 270786
rect 118025 270752 118297 270786
rect 118425 270752 118697 270786
rect 118825 270752 118841 270786
rect 115648 270715 118841 270752
rect 115648 270714 115700 270715
rect 114050 270673 114542 270693
rect 114050 270576 114086 270673
rect 114501 270576 114542 270673
rect 114050 270545 114542 270576
rect 114364 270296 114537 270545
rect 118418 270296 118934 270326
rect 112560 270262 112576 270296
rect 112704 270262 112976 270296
rect 113104 270262 113376 270296
rect 113504 270262 113776 270296
rect 113904 270262 114176 270296
rect 114304 270262 114576 270296
rect 114704 270262 114976 270296
rect 115104 270262 115376 270296
rect 115504 270262 115776 270296
rect 115904 270262 116176 270296
rect 116304 270262 116576 270296
rect 116704 270262 116976 270296
rect 117104 270262 117376 270296
rect 117504 270262 117776 270296
rect 117904 270262 118176 270296
rect 118304 270262 118576 270296
rect 118704 270288 118934 270296
rect 118704 270262 118720 270288
rect 112514 270212 112548 270228
rect 112514 269120 112548 269136
rect 112732 270212 112766 270228
rect 112732 269120 112766 269136
rect 112914 270212 112948 270228
rect 112914 269120 112948 269136
rect 113132 270212 113166 270228
rect 113132 269120 113166 269136
rect 113314 270212 113348 270228
rect 113314 269120 113348 269136
rect 113532 270212 113566 270228
rect 113532 269120 113566 269136
rect 113714 270212 113748 270228
rect 113714 269120 113748 269136
rect 113932 270212 113966 270228
rect 113932 269120 113966 269136
rect 114114 270212 114148 270228
rect 114114 269120 114148 269136
rect 114332 270212 114366 270228
rect 114332 269120 114366 269136
rect 114514 270212 114548 270228
rect 114514 269120 114548 269136
rect 114732 270212 114766 270228
rect 114732 269120 114766 269136
rect 114914 270212 114948 270228
rect 114914 269120 114948 269136
rect 115132 270212 115166 270228
rect 115132 269120 115166 269136
rect 115314 270212 115348 270228
rect 115314 269120 115348 269136
rect 115532 270212 115566 270228
rect 115532 269120 115566 269136
rect 115714 270212 115748 270228
rect 115714 269120 115748 269136
rect 115932 270212 115966 270228
rect 115932 269120 115966 269136
rect 116114 270212 116148 270228
rect 116114 269120 116148 269136
rect 116332 270212 116366 270228
rect 116332 269120 116366 269136
rect 116514 270212 116548 270228
rect 116514 269120 116548 269136
rect 116732 270212 116766 270228
rect 116732 269120 116766 269136
rect 116914 270212 116948 270228
rect 116914 269120 116948 269136
rect 117132 270212 117166 270228
rect 117132 269120 117166 269136
rect 117314 270212 117348 270228
rect 117314 269120 117348 269136
rect 117532 270212 117566 270228
rect 117532 269120 117566 269136
rect 117714 270212 117748 270228
rect 117714 269120 117748 269136
rect 117932 270212 117966 270228
rect 117932 269120 117966 269136
rect 118114 270212 118148 270228
rect 118114 269120 118148 269136
rect 118332 270212 118366 270228
rect 118332 269120 118366 269136
rect 118514 270212 118548 270228
rect 118514 269120 118548 269136
rect 118732 270212 118766 270228
rect 118732 269120 118766 269136
rect 112560 269052 112576 269086
rect 112704 269052 112976 269086
rect 113104 269052 113376 269086
rect 113504 269052 113776 269086
rect 113904 269052 114176 269086
rect 114304 269052 114576 269086
rect 114704 269052 114976 269086
rect 115104 269052 115376 269086
rect 115504 269052 115776 269086
rect 115904 269052 116176 269086
rect 116304 269052 116576 269086
rect 116704 269052 116976 269086
rect 117104 269052 117376 269086
rect 117504 269052 117776 269086
rect 117904 269052 118176 269086
rect 118304 269052 118576 269086
rect 118704 269055 118720 269086
rect 118882 269055 118934 270288
rect 118704 269052 118934 269055
rect 118416 269017 118934 269052
rect 114230 268883 117626 268907
rect 114230 268826 114322 268883
rect 117498 268826 117626 268883
rect 112069 268702 112160 268826
rect 118949 268702 119021 268826
rect 112069 268675 119021 268702
rect 119151 272179 119158 272249
rect 120104 281012 120227 281067
rect 125148 281012 125658 281165
rect 125047 280856 125658 281012
rect 120237 280779 120297 280813
rect 121668 280800 121728 280813
rect 121668 280779 121960 280800
rect 120237 280753 121960 280779
rect 120271 280718 121694 280753
rect 120271 280684 120445 280718
rect 120813 280713 121145 280718
rect 120813 280684 120875 280713
rect 120271 280641 120429 280684
rect 120829 280641 120875 280684
rect 120271 280625 120417 280641
rect 120271 280549 120383 280625
rect 120271 280533 120417 280549
rect 120841 280625 120875 280641
rect 120841 280533 120875 280549
rect 121083 280684 121145 280713
rect 121513 280684 121694 280718
rect 121083 280641 121129 280684
rect 121529 280641 121694 280684
rect 121083 280625 121117 280641
rect 121083 280533 121117 280549
rect 121541 280625 121694 280641
rect 121575 280549 121694 280625
rect 121541 280545 121694 280549
rect 121541 280533 121575 280545
rect 120271 280257 120395 280533
rect 120429 280456 120445 280490
rect 120813 280456 120829 280490
rect 121129 280456 121145 280490
rect 121513 280456 121529 280490
rect 120429 280300 120445 280334
rect 120813 280300 120829 280334
rect 121129 280300 121145 280334
rect 121513 280300 121529 280334
rect 120271 280241 120417 280257
rect 120271 279765 120383 280241
rect 120271 279749 120417 279765
rect 120841 280241 120875 280257
rect 120841 279749 120875 279765
rect 121083 280241 121117 280257
rect 121083 279749 121117 279765
rect 121541 280241 121575 280257
rect 121541 279749 121575 279765
rect 120271 279473 120395 279749
rect 120429 279672 120445 279706
rect 120813 279672 120829 279706
rect 121129 279672 121145 279706
rect 121513 279672 121529 279706
rect 120429 279516 120445 279550
rect 120813 279516 120829 279550
rect 121129 279516 121145 279550
rect 121513 279516 121529 279550
rect 120271 279457 120417 279473
rect 120271 278981 120383 279457
rect 120271 278965 120417 278981
rect 120841 279457 120875 279473
rect 120841 278965 120875 278981
rect 121083 279457 121117 279473
rect 121083 278965 121117 278981
rect 121541 279457 121575 279473
rect 121541 278965 121575 278981
rect 120271 278689 120395 278965
rect 120429 278888 120445 278922
rect 120813 278888 120829 278922
rect 121129 278888 121145 278922
rect 121513 278888 121529 278922
rect 120429 278732 120445 278766
rect 120813 278732 120829 278766
rect 121129 278732 121145 278766
rect 121513 278732 121529 278766
rect 120271 278673 120417 278689
rect 120271 278197 120383 278673
rect 120271 278181 120417 278197
rect 120841 278673 120875 278689
rect 120841 278181 120875 278197
rect 121083 278673 121117 278689
rect 121083 278181 121117 278197
rect 121541 278673 121575 278689
rect 121541 278181 121575 278197
rect 120271 277905 120395 278181
rect 120429 278104 120445 278138
rect 120813 278104 120829 278138
rect 121129 278104 121145 278138
rect 121513 278104 121529 278138
rect 120429 277948 120445 277982
rect 120813 277948 120829 277982
rect 121129 277948 121145 277982
rect 121513 277948 121529 277982
rect 120271 277889 120417 277905
rect 120271 277413 120383 277889
rect 120271 277397 120417 277413
rect 120841 277889 120875 277905
rect 120841 277397 120875 277413
rect 121083 277889 121117 277905
rect 121083 277397 121117 277413
rect 121541 277889 121575 277905
rect 121541 277397 121575 277413
rect 120271 277121 120395 277397
rect 120429 277320 120445 277354
rect 120813 277320 120829 277354
rect 121129 277320 121145 277354
rect 121513 277320 121529 277354
rect 120429 277164 120445 277198
rect 120813 277164 120829 277198
rect 121129 277164 121145 277198
rect 121513 277164 121529 277198
rect 120271 277105 120417 277121
rect 120271 276629 120383 277105
rect 120271 276613 120417 276629
rect 120841 277105 120875 277121
rect 120841 276613 120875 276629
rect 121083 277105 121117 277121
rect 121083 276613 121117 276629
rect 121541 277105 121575 277121
rect 121541 276613 121575 276629
rect 120271 276337 120395 276613
rect 120429 276536 120445 276570
rect 120813 276536 120829 276570
rect 121129 276536 121145 276570
rect 121513 276536 121529 276570
rect 120429 276380 120445 276414
rect 120813 276380 120829 276414
rect 121129 276380 121145 276414
rect 121513 276380 121529 276414
rect 120271 276321 120417 276337
rect 120271 275845 120383 276321
rect 120271 275829 120417 275845
rect 120841 276321 120875 276337
rect 121083 276321 121117 276337
rect 120875 276118 121083 276139
rect 120875 276054 120958 276118
rect 121014 276054 121083 276118
rect 120875 276032 121083 276054
rect 120841 275829 120875 275845
rect 121083 275829 121117 275845
rect 121541 276321 121575 276337
rect 121541 275829 121575 275845
rect 120271 275553 120395 275829
rect 120429 275752 120445 275786
rect 120813 275752 120829 275786
rect 121129 275752 121145 275786
rect 121513 275752 121529 275786
rect 120429 275596 120445 275630
rect 120813 275596 120829 275630
rect 121129 275596 121145 275630
rect 121513 275596 121529 275630
rect 120271 275537 120417 275553
rect 120271 275061 120383 275537
rect 120271 275045 120417 275061
rect 120841 275537 120875 275553
rect 121083 275537 121117 275553
rect 120875 275246 121083 275353
rect 120841 275045 120875 275061
rect 120271 274769 120395 275045
rect 120429 274968 120445 275002
rect 120813 274968 120829 275002
rect 120429 274812 120445 274846
rect 120813 274812 120829 274846
rect 120271 274753 120417 274769
rect 120271 274277 120383 274753
rect 120271 274261 120417 274277
rect 120841 274753 120875 274769
rect 120943 274579 121039 275246
rect 121083 275045 121117 275061
rect 121541 275537 121575 275553
rect 121541 275045 121575 275061
rect 121129 274968 121145 275002
rect 121513 274968 121529 275002
rect 121129 274812 121145 274846
rect 121513 274812 121529 274846
rect 121083 274753 121117 274769
rect 120875 274472 121083 274579
rect 120841 274261 120875 274277
rect 121083 274261 121117 274277
rect 121541 274753 121575 274769
rect 121541 274261 121575 274277
rect 120271 273985 120395 274261
rect 120429 274184 120445 274218
rect 120813 274184 120829 274218
rect 121129 274184 121145 274218
rect 121513 274184 121529 274218
rect 120429 274028 120445 274062
rect 120813 274028 120829 274062
rect 121129 274028 121145 274062
rect 121513 274028 121529 274062
rect 120271 273969 120417 273985
rect 120271 273493 120383 273969
rect 120271 273477 120417 273493
rect 120841 273969 120875 273985
rect 121083 273969 121117 273985
rect 120875 273756 121083 273778
rect 120875 273692 120961 273756
rect 121017 273692 121083 273756
rect 120875 273671 121083 273692
rect 120841 273477 120875 273493
rect 121083 273477 121117 273493
rect 121541 273969 121575 273985
rect 121541 273477 121575 273493
rect 120271 273201 120395 273477
rect 120429 273400 120445 273434
rect 120813 273400 120829 273434
rect 121129 273400 121145 273434
rect 121513 273400 121529 273434
rect 120429 273244 120445 273278
rect 120813 273244 120829 273278
rect 121129 273244 121145 273278
rect 121513 273244 121529 273278
rect 120271 273185 120417 273201
rect 120271 272709 120383 273185
rect 120271 272693 120417 272709
rect 120841 273185 120875 273201
rect 120841 272693 120875 272709
rect 121083 273185 121117 273201
rect 121083 272693 121117 272709
rect 121541 273185 121575 273201
rect 121541 272693 121575 272709
rect 120271 272417 120395 272693
rect 120429 272616 120445 272650
rect 120813 272616 120829 272650
rect 121129 272616 121145 272650
rect 121513 272616 121529 272650
rect 120429 272460 120445 272494
rect 120813 272460 120829 272494
rect 121129 272460 121145 272494
rect 121513 272460 121529 272494
rect 120271 272401 120417 272417
rect 120271 271925 120383 272401
rect 120271 271909 120417 271925
rect 120841 272401 120875 272417
rect 120841 271909 120875 271925
rect 121083 272401 121117 272417
rect 121083 271909 121117 271925
rect 121541 272401 121575 272417
rect 121541 271909 121575 271925
rect 120271 271633 120395 271909
rect 120429 271832 120445 271866
rect 120813 271832 120829 271866
rect 121129 271832 121145 271866
rect 121513 271832 121529 271866
rect 120429 271676 120445 271710
rect 120813 271676 120829 271710
rect 121129 271676 121145 271710
rect 121513 271676 121529 271710
rect 120271 271617 120417 271633
rect 120271 271141 120383 271617
rect 120271 271125 120417 271141
rect 120841 271617 120875 271633
rect 120841 271125 120875 271141
rect 121083 271617 121117 271633
rect 121083 271125 121117 271141
rect 121541 271617 121575 271633
rect 121541 271125 121575 271141
rect 120271 270849 120395 271125
rect 120429 271048 120445 271082
rect 120813 271048 120829 271082
rect 121129 271048 121145 271082
rect 121513 271048 121529 271082
rect 120429 270892 120445 270926
rect 120813 270892 120829 270926
rect 121129 270892 121145 270926
rect 121513 270892 121529 270926
rect 120271 270833 120417 270849
rect 120271 270357 120383 270833
rect 120271 270341 120417 270357
rect 120841 270833 120875 270849
rect 120841 270341 120875 270357
rect 121083 270833 121117 270849
rect 121083 270341 121117 270357
rect 121541 270833 121575 270849
rect 121541 270341 121575 270357
rect 120271 270065 120395 270341
rect 120429 270264 120445 270298
rect 120813 270264 120829 270298
rect 121129 270264 121145 270298
rect 121513 270264 121529 270298
rect 120429 270108 120445 270142
rect 120813 270108 120829 270142
rect 121129 270108 121145 270142
rect 121513 270108 121529 270142
rect 120271 270049 120417 270065
rect 120271 269573 120383 270049
rect 120271 269557 120417 269573
rect 120841 270049 120875 270065
rect 120841 269557 120875 269573
rect 121083 270049 121117 270065
rect 121083 269557 121117 269573
rect 121541 270049 121575 270065
rect 121541 269557 121575 269573
rect 120271 269281 120395 269557
rect 120429 269480 120445 269514
rect 120813 269480 120829 269514
rect 121129 269480 121145 269514
rect 121513 269480 121529 269514
rect 120429 269324 120445 269358
rect 120813 269324 120829 269358
rect 121129 269324 121145 269358
rect 121513 269324 121529 269358
rect 120271 269265 120417 269281
rect 120271 269189 120383 269265
rect 120271 269173 120417 269189
rect 120841 269265 120875 269281
rect 120841 269173 120875 269189
rect 120271 269130 120429 269173
rect 120829 269130 120875 269173
rect 120271 269096 120445 269130
rect 120813 269114 120875 269130
rect 121083 269265 121117 269281
rect 121083 269173 121117 269189
rect 121541 269265 121575 269281
rect 121541 269173 121575 269189
rect 121083 269130 121129 269173
rect 121529 269130 121575 269173
rect 121083 269114 121145 269130
rect 120813 269096 121145 269114
rect 121513 269114 121575 269130
rect 121513 269096 121694 269114
rect 120271 269038 121694 269096
rect 121728 279988 121960 280753
rect 122178 280574 122238 280608
rect 123578 280574 123638 280608
rect 122178 280548 122212 280574
rect 121728 279887 122178 279988
rect 123604 280548 123638 280574
rect 122356 280470 122372 280504
rect 122740 280470 122756 280504
rect 123056 280470 123072 280504
rect 123440 280470 123456 280504
rect 122212 280411 122344 280427
rect 122212 279935 122310 280411
rect 122212 279919 122344 279935
rect 122768 280411 122802 280427
rect 122768 279919 122802 279935
rect 123010 280411 123044 280427
rect 123010 279919 123044 279935
rect 123468 280411 123502 280427
rect 123468 279919 123502 279935
rect 121728 279275 121849 279887
rect 122212 279643 122310 279919
rect 122356 279842 122372 279876
rect 122740 279842 122756 279876
rect 123056 279842 123072 279876
rect 123440 279842 123456 279876
rect 122356 279686 122372 279720
rect 122740 279686 122756 279720
rect 123056 279686 123072 279720
rect 123440 279686 123456 279720
rect 122212 279627 122344 279643
rect 121728 279026 122178 279275
rect 122212 279151 122310 279627
rect 122212 279135 122344 279151
rect 122768 279627 122802 279643
rect 122768 279135 122802 279151
rect 123010 279627 123044 279643
rect 123010 279135 123044 279151
rect 123468 279627 123502 279643
rect 123468 279135 123502 279151
rect 122356 279058 122372 279092
rect 122740 279058 122756 279092
rect 123056 279058 123072 279092
rect 123440 279058 123456 279092
rect 121728 279000 122212 279026
rect 123604 279000 123638 279026
rect 121728 278966 122238 279000
rect 123578 278966 123638 279000
rect 121728 278870 123358 278966
rect 121728 273057 121809 278870
rect 122027 278619 122144 278635
rect 122022 276038 122027 276225
rect 122260 278482 123358 278870
rect 122254 278448 122314 278482
rect 124310 278448 124370 278482
rect 122254 278422 122374 278448
rect 122288 278270 122374 278422
rect 124336 278422 124370 278448
rect 122414 278313 122430 278347
rect 123274 278313 123290 278347
rect 122288 278254 122402 278270
rect 122288 277804 122368 278254
rect 122288 277788 122402 277804
rect 123302 278254 123336 278270
rect 123336 278161 124210 278193
rect 123336 278154 123672 278161
rect 123302 277788 123336 277804
rect 122288 277504 122374 277788
rect 122414 277711 122430 277745
rect 123274 277711 123290 277745
rect 122416 277547 122432 277581
rect 123200 277547 123216 277581
rect 122288 277488 122404 277504
rect 122288 277412 122370 277488
rect 122288 277396 122404 277412
rect 123228 277488 123262 277504
rect 123228 277396 123262 277412
rect 122288 277247 122374 277396
rect 122416 277319 122432 277353
rect 123200 277319 123216 277353
rect 123494 277330 123535 278154
rect 123656 278127 123672 278154
rect 124194 278127 124210 278161
rect 123610 278068 123644 278084
rect 123610 277390 123644 277406
rect 124222 278068 124256 278084
rect 124222 277390 124256 277406
rect 123656 277330 123672 277347
rect 123494 277313 123672 277330
rect 124194 277313 124210 277347
rect 123494 277290 124210 277313
rect 122254 277221 122374 277247
rect 124336 277221 124370 277247
rect 122254 277187 122314 277221
rect 124310 277187 124370 277221
rect 123686 277034 123945 277076
rect 123686 276881 123736 277034
rect 123913 276881 123945 277034
rect 123686 276851 123945 276881
rect 122278 276817 122374 276851
rect 123896 276817 123992 276851
rect 122278 276755 123860 276817
rect 122312 276749 123860 276755
rect 122312 276715 122454 276749
rect 123816 276740 123860 276749
rect 123958 276755 123992 276817
rect 123816 276715 123832 276740
rect 122312 276656 122426 276715
rect 122312 276504 122392 276656
rect 122312 276445 122426 276504
rect 123844 276656 123878 276672
rect 123844 276488 123878 276504
rect 122312 276411 122454 276445
rect 123816 276419 123832 276445
rect 123816 276411 123862 276419
rect 122312 276405 123862 276411
rect 122278 276343 123862 276405
rect 123958 276343 123992 276405
rect 122278 276309 122374 276343
rect 123896 276309 123992 276343
rect 124173 276382 125047 276742
rect 122144 276212 122552 276225
rect 124173 276212 124291 276382
rect 122144 276131 122500 276212
rect 122404 276097 122500 276131
rect 124297 276097 124313 276212
rect 122404 276060 122552 276097
rect 122144 276038 122552 276060
rect 124445 276083 124567 276110
rect 122144 276035 122427 276038
rect 124445 275982 124465 276083
rect 124549 275982 124567 276083
rect 124445 275971 124567 275982
rect 122283 275937 122379 275971
rect 124861 275937 124957 275971
rect 122283 275875 122317 275937
rect 124923 275875 124957 275937
rect 122462 275823 122478 275857
rect 122854 275823 122870 275857
rect 123098 275823 123114 275857
rect 123490 275823 123506 275857
rect 123734 275823 123750 275857
rect 124126 275823 124142 275857
rect 124370 275823 124386 275857
rect 124762 275823 124778 275857
rect 122385 275795 122419 275811
rect 122385 275711 122419 275727
rect 122913 275795 122947 275811
rect 122913 275711 122947 275727
rect 123021 275795 123055 275811
rect 123021 275711 123055 275727
rect 123549 275795 123583 275811
rect 123549 275711 123583 275727
rect 123657 275795 123691 275811
rect 123657 275711 123691 275727
rect 124185 275795 124219 275811
rect 124185 275711 124219 275727
rect 124293 275795 124327 275811
rect 124293 275711 124327 275727
rect 124821 275795 124855 275811
rect 124821 275711 124855 275727
rect 122283 275585 122317 275647
rect 122462 275665 122478 275699
rect 122854 275665 122870 275699
rect 122462 275585 122870 275665
rect 123098 275665 123114 275699
rect 123490 275665 123506 275699
rect 123098 275585 123506 275665
rect 123734 275665 123750 275699
rect 124126 275665 124142 275699
rect 123734 275585 124142 275665
rect 124370 275665 124386 275699
rect 124762 275665 124778 275699
rect 124370 275585 124778 275665
rect 124923 275585 124957 275647
rect 122283 275551 122379 275585
rect 124861 275551 124957 275585
rect 122027 275515 122144 275531
rect 123246 275431 123421 275551
rect 123213 275386 123457 275431
rect 123213 275173 123245 275386
rect 123426 275173 123457 275386
rect 123213 275140 123457 275173
rect 122792 275002 122888 275036
rect 124016 275002 124112 275036
rect 122792 274940 122826 275002
rect 124078 274940 124112 275002
rect 122952 274900 122968 274934
rect 123936 274900 123952 274934
rect 122906 274850 122940 274866
rect 122906 274658 122940 274674
rect 123964 274850 123998 274866
rect 123998 274715 124078 274816
rect 123964 274658 123998 274674
rect 122952 274590 122968 274624
rect 123936 274590 123952 274624
rect 122792 274562 122826 274584
rect 122060 274486 122084 274562
rect 122714 274522 122826 274562
rect 124078 274537 124112 274584
rect 124202 274537 124218 274582
rect 124078 274522 124218 274537
rect 122714 274488 122888 274522
rect 124016 274488 124218 274522
rect 124824 274555 124840 274582
rect 124824 274488 125047 274555
rect 122714 274486 122730 274488
rect 122060 274354 122253 274486
rect 122523 274354 122558 274392
rect 122061 274350 122558 274354
rect 122061 274316 122293 274350
rect 122461 274316 122558 274350
rect 122693 274316 122709 274350
rect 122877 274316 122893 274350
rect 122061 274296 122558 274316
rect 122061 274282 122062 274296
rect 122150 274282 122558 274296
rect 122939 274282 122974 274488
rect 123497 274445 123670 274452
rect 123497 274437 123527 274445
rect 123354 274408 123527 274437
rect 123647 274437 123670 274445
rect 123647 274408 123806 274437
rect 123354 274399 123806 274408
rect 123354 274387 123390 274399
rect 123109 274316 123125 274350
rect 123293 274316 123309 274350
rect 123355 274282 123390 274387
rect 123525 274316 123541 274350
rect 123709 274316 123725 274350
rect 123771 274282 123806 274399
rect 123941 274316 123957 274350
rect 124125 274316 124141 274350
rect 124187 274282 124222 274488
rect 124603 274354 124638 274392
rect 124726 274354 125047 274488
rect 122150 274266 122265 274282
rect 122150 273790 122231 274266
rect 122150 273774 122265 273790
rect 122489 274266 122558 274282
rect 122523 273790 122558 274266
rect 122489 273774 122558 273790
rect 122647 274266 122681 274282
rect 122647 273774 122681 273790
rect 122905 274266 122974 274282
rect 122939 273790 122974 274266
rect 122905 273774 122974 273790
rect 123063 274266 123097 274282
rect 123063 273774 123097 273790
rect 123321 274266 123390 274282
rect 123355 273790 123390 274266
rect 123321 273774 123390 273790
rect 123479 274266 123513 274282
rect 123479 273774 123513 273790
rect 123737 274266 123806 274282
rect 123771 273790 123806 274266
rect 123737 273774 123806 273790
rect 123895 274266 123929 274282
rect 123895 273774 123929 273790
rect 124153 274266 124222 274282
rect 124187 273790 124222 274266
rect 124153 273774 124222 273790
rect 124311 274350 125047 274354
rect 124311 274316 124373 274350
rect 124541 274316 125047 274350
rect 124311 274312 125047 274316
rect 124311 274282 124726 274312
rect 124311 274266 124345 274282
rect 124311 273774 124345 273790
rect 124569 274266 124726 274282
rect 124603 273790 124726 274266
rect 124569 273774 124726 273790
rect 122150 273740 122558 273774
rect 124311 273740 124726 273774
rect 122150 273706 122293 273740
rect 122461 273706 122558 273740
rect 122693 273706 122709 273740
rect 122877 273706 122893 273740
rect 123109 273706 123125 273740
rect 123293 273706 123309 273740
rect 123525 273706 123541 273740
rect 123709 273706 123725 273740
rect 123941 273706 123957 273740
rect 124125 273706 124141 273740
rect 124311 273706 124373 273740
rect 124541 273706 124726 273740
rect 122150 273702 122558 273706
rect 124311 273702 124726 273706
rect 122150 273621 122253 273702
rect 122062 273618 122253 273621
rect 124610 273637 124726 273702
rect 124814 273637 125047 274312
rect 124610 273618 125047 273637
rect 122062 273545 122217 273618
rect 124615 273545 125047 273618
rect 121728 272998 123538 273057
rect 121728 272964 121980 272998
rect 123494 272964 123554 272998
rect 121728 272954 123554 272964
rect 121728 272938 121954 272954
rect 121728 269054 121920 272938
rect 122079 272894 122571 272954
rect 122079 272860 122141 272894
rect 122509 272860 122571 272894
rect 122079 272801 122125 272860
rect 122113 272725 122125 272801
rect 122079 272666 122125 272725
rect 122525 272801 122571 272860
rect 122525 272725 122537 272801
rect 122525 272666 122571 272725
rect 122079 272632 122141 272666
rect 122509 272632 122571 272666
rect 122779 272894 123271 272954
rect 122779 272860 122841 272894
rect 123209 272860 123271 272894
rect 122779 272801 122825 272860
rect 122813 272725 122825 272801
rect 122779 272666 122825 272725
rect 123225 272801 123271 272860
rect 123225 272725 123237 272801
rect 123225 272666 123271 272725
rect 122779 272632 122841 272666
rect 123209 272632 123271 272666
rect 123520 272938 123554 272954
rect 123333 272626 123462 272656
rect 123333 272510 123355 272626
rect 122125 272476 122141 272510
rect 122509 272476 122525 272510
rect 122825 272476 122841 272510
rect 123209 272476 123355 272510
rect 123333 272446 123355 272476
rect 123444 272446 123462 272626
rect 122079 272417 122113 272433
rect 121954 272123 122079 272248
rect 122079 271925 122113 271941
rect 122537 272417 122571 272433
rect 122779 272417 122813 272433
rect 122571 272214 122779 272235
rect 122571 272150 122654 272214
rect 122710 272150 122779 272214
rect 122571 272128 122779 272150
rect 122537 271925 122571 271941
rect 122779 271925 122813 271941
rect 123237 272417 123271 272433
rect 123237 271925 123271 271941
rect 123333 272427 123462 272446
rect 123333 271882 123367 272427
rect 122125 271848 122141 271882
rect 122509 271848 122525 271882
rect 122825 271848 122841 271882
rect 123209 271848 123367 271882
rect 122125 271692 122141 271726
rect 122509 271692 122525 271726
rect 122825 271692 122841 271726
rect 123209 271692 123225 271726
rect 122079 271633 122113 271649
rect 121954 271331 122079 271456
rect 122079 271141 122113 271157
rect 122537 271633 122571 271649
rect 122779 271633 122813 271649
rect 122571 271342 122779 271449
rect 122537 271141 122571 271157
rect 122125 271064 122141 271098
rect 122509 271064 122525 271098
rect 122125 270908 122141 270942
rect 122509 270908 122525 270942
rect 122079 270849 122113 270865
rect 121954 270547 122079 270672
rect 122079 270357 122113 270373
rect 122537 270849 122571 270865
rect 122639 270675 122735 271342
rect 122779 271141 122813 271157
rect 123237 271633 123271 271649
rect 123237 271141 123271 271157
rect 122825 271064 122841 271098
rect 123209 271064 123225 271098
rect 122825 270908 122841 270942
rect 123209 270908 123225 270942
rect 122779 270849 122813 270865
rect 122571 270568 122779 270675
rect 122537 270357 122571 270373
rect 122779 270357 122813 270373
rect 123237 270849 123271 270865
rect 123237 270357 123271 270373
rect 122125 270280 122141 270314
rect 122509 270280 122525 270314
rect 122825 270280 122841 270314
rect 123209 270280 123225 270314
rect 122125 270124 122141 270158
rect 122509 270124 122525 270158
rect 122825 270124 122841 270158
rect 123209 270124 123351 270158
rect 122079 270065 122113 270081
rect 121954 269757 122079 269882
rect 122079 269573 122113 269589
rect 122537 270065 122571 270081
rect 122779 270065 122813 270081
rect 122571 269852 122779 269874
rect 122571 269788 122657 269852
rect 122713 269788 122779 269852
rect 122571 269767 122779 269788
rect 122537 269573 122571 269589
rect 122779 269573 122813 269589
rect 123237 270065 123271 270081
rect 123237 269573 123271 269589
rect 123317 269530 123351 270124
rect 122125 269496 122141 269530
rect 122509 269496 122525 269530
rect 122825 269496 122841 269530
rect 123209 269496 123351 269530
rect 122079 269340 122141 269374
rect 122509 269340 122571 269374
rect 122079 269281 122125 269340
rect 122113 269205 122125 269281
rect 122079 269146 122125 269205
rect 122525 269281 122571 269340
rect 122525 269205 122537 269281
rect 122525 269146 122571 269205
rect 122079 269112 122141 269146
rect 122509 269112 122571 269146
rect 122079 269066 122571 269112
rect 122779 269340 122841 269374
rect 123209 269340 123271 269374
rect 122779 269281 122825 269340
rect 122813 269205 122825 269281
rect 122779 269146 122825 269205
rect 123225 269281 123271 269340
rect 123225 269205 123237 269281
rect 123225 269146 123271 269205
rect 122779 269112 122841 269146
rect 123209 269112 123271 269146
rect 122779 269066 123271 269112
rect 121954 269054 123520 269066
rect 121728 269038 123554 269054
rect 120237 269028 123554 269038
rect 120237 269012 121980 269028
rect 120237 268978 120297 269012
rect 121668 268994 121980 269012
rect 123494 268994 123554 269028
rect 123827 272777 124279 273545
rect 123827 272689 124051 272777
rect 124726 272770 124768 272777
rect 124726 272717 125047 272770
rect 124726 272689 124811 272717
rect 123827 272598 124029 272689
rect 123827 269356 123978 272598
rect 124116 272601 124188 272689
rect 124696 272601 124811 272689
rect 124116 272566 124811 272601
rect 124116 272532 124204 272566
rect 124680 272532 124768 272566
rect 124116 272504 124188 272532
rect 124116 272336 124120 272504
rect 124154 272336 124188 272504
rect 124116 272308 124188 272336
rect 124696 272504 124768 272532
rect 124696 272336 124730 272504
rect 124764 272336 124768 272504
rect 124696 272308 124768 272336
rect 124116 272274 124204 272308
rect 124680 272274 124768 272308
rect 124188 272150 124811 272185
rect 124188 272116 124204 272150
rect 124680 272116 124696 272150
rect 124084 272088 124154 272104
rect 124084 271920 124120 272088
rect 124084 271904 124154 271920
rect 124730 272088 124764 272104
rect 124730 271904 124764 271920
rect 124084 271688 124120 271904
rect 124188 271858 124204 271892
rect 124680 271858 124696 271892
rect 124188 271734 124811 271769
rect 124188 271700 124204 271734
rect 124680 271700 124696 271734
rect 124084 271672 124154 271688
rect 124084 271504 124120 271672
rect 124084 271488 124154 271504
rect 124730 271672 124764 271688
rect 124730 271488 124764 271504
rect 124084 271272 124120 271488
rect 124188 271442 124204 271476
rect 124680 271442 124696 271476
rect 124188 271318 124811 271353
rect 124188 271284 124204 271318
rect 124680 271284 124696 271318
rect 124084 271256 124154 271272
rect 124084 271088 124120 271256
rect 124084 271072 124154 271088
rect 124730 271256 124764 271272
rect 124730 271072 124764 271088
rect 124084 270856 124120 271072
rect 124188 271026 124204 271060
rect 124680 271026 124696 271060
rect 124188 270902 124811 270937
rect 124188 270868 124204 270902
rect 124680 270868 124696 270902
rect 124084 270840 124154 270856
rect 124084 270672 124120 270840
rect 124084 270656 124154 270672
rect 124730 270840 124764 270856
rect 124730 270656 124764 270672
rect 124084 270440 124120 270656
rect 124188 270610 124204 270644
rect 124680 270610 124696 270644
rect 124188 270486 124811 270521
rect 124188 270452 124204 270486
rect 124680 270452 124696 270486
rect 124084 270424 124154 270440
rect 124084 270256 124120 270424
rect 124084 270240 124154 270256
rect 124730 270424 124764 270440
rect 124730 270240 124764 270256
rect 124084 270024 124120 270240
rect 124188 270194 124204 270228
rect 124680 270194 124696 270228
rect 124188 270070 124811 270105
rect 124188 270036 124204 270070
rect 124680 270036 124696 270070
rect 124084 270008 124154 270024
rect 124084 269840 124120 270008
rect 124084 269824 124154 269840
rect 124730 270008 124764 270024
rect 124730 269824 124764 269840
rect 124188 269778 124204 269812
rect 124680 269778 124696 269812
rect 123827 269281 124029 269356
rect 124116 269654 124811 269689
rect 124116 269620 124204 269654
rect 124680 269620 124811 269654
rect 124116 269592 124188 269620
rect 124116 269424 124120 269592
rect 124154 269424 124188 269592
rect 124116 269396 124188 269424
rect 124696 269592 124811 269620
rect 124696 269424 124730 269592
rect 124764 269424 124811 269592
rect 124696 269396 124811 269424
rect 124116 269362 124204 269396
rect 124680 269362 124811 269396
rect 124116 269281 124188 269362
rect 124696 269291 124811 269362
rect 124880 272580 125047 272717
rect 124880 269291 125047 269668
rect 124696 269281 125047 269291
rect 123827 269193 124035 269281
rect 124710 269193 125047 269281
rect 121668 268978 123550 268994
rect 120307 268946 123550 268978
rect 121789 268938 123550 268946
rect 123827 268990 125047 269193
rect 125171 275523 125658 280856
rect 125171 275158 128452 275523
rect 125171 268990 125790 275158
rect 123827 268861 125790 268990
rect 120104 268778 120254 268861
rect 119938 268708 120254 268778
rect 125175 268708 125790 268861
rect 111939 268659 119151 268675
rect 112005 268607 119104 268659
rect 123847 268607 125790 268708
rect 105957 268342 125790 268607
rect 128055 268342 128452 275158
rect 105957 268022 128452 268342
rect 105957 268007 125658 268022
<< viali >>
rect 106373 280851 106473 280885
rect 106773 280851 106873 280885
rect 107173 280851 107273 280885
rect 107573 280851 107673 280885
rect 107973 280851 108073 280885
rect 108373 280851 108473 280885
rect 108773 280851 108873 280885
rect 109173 280851 109273 280885
rect 109573 280851 109673 280885
rect 109973 280851 110073 280885
rect 106311 279805 106345 280801
rect 106501 279805 106535 280801
rect 106711 279805 106745 280801
rect 106901 279805 106935 280801
rect 107111 279805 107145 280801
rect 107301 279805 107335 280801
rect 107511 279805 107545 280801
rect 107701 279805 107735 280801
rect 107911 279805 107945 280801
rect 108101 279805 108135 280801
rect 108311 279805 108345 280801
rect 108501 279805 108535 280801
rect 108711 279805 108745 280801
rect 108901 279805 108935 280801
rect 109111 279805 109145 280801
rect 109301 279805 109335 280801
rect 109511 279805 109545 280801
rect 109701 279805 109735 280801
rect 109911 279805 109945 280801
rect 110101 279805 110135 280801
rect 106373 279721 106473 279755
rect 106773 279721 106873 279755
rect 107173 279721 107273 279755
rect 107573 279721 107673 279755
rect 107973 279721 108073 279755
rect 108373 279721 108473 279755
rect 108773 279721 108873 279755
rect 109173 279721 109273 279755
rect 109573 279721 109673 279755
rect 109973 279721 110073 279755
rect 106380 279023 107570 279057
rect 106287 278773 106321 278995
rect 107629 278773 107663 278995
rect 106380 278711 107570 278745
rect 106380 278423 107570 278457
rect 106287 278173 106321 278395
rect 107629 278173 107663 278395
rect 106380 278111 107570 278145
rect 106941 277984 107098 278068
rect 106941 277950 107098 277984
rect 106941 277789 107098 277950
rect 106503 277176 107513 277210
rect 106410 277106 106444 277148
rect 107572 277106 107606 277148
rect 106503 277044 107513 277078
rect 109793 279049 110047 279083
rect 109731 277985 109765 278999
rect 110075 277985 110109 278999
rect 109793 277901 110047 277935
rect 109793 277793 110047 277827
rect 109731 276729 109765 277743
rect 110075 276729 110109 277743
rect 109793 276645 110047 276679
rect 106375 274853 106549 276290
rect 106963 275725 107117 275759
rect 107463 275725 107617 275759
rect 107963 275725 108117 275759
rect 108463 275725 108617 275759
rect 108963 275725 109117 275759
rect 109463 275725 109617 275759
rect 106870 274951 106904 275697
rect 107176 274951 107210 275697
rect 107370 274951 107404 275697
rect 107676 274951 107710 275697
rect 107870 274951 107904 275697
rect 108176 274951 108210 275697
rect 108370 274951 108404 275697
rect 108676 274951 108710 275697
rect 108870 274951 108904 275697
rect 109176 274951 109210 275697
rect 109370 274951 109404 275697
rect 109676 274951 109710 275697
rect 106963 274889 107117 274923
rect 107463 274889 107617 274923
rect 107963 274889 108117 274923
rect 108463 274889 108617 274923
rect 108963 274889 109117 274923
rect 109463 274889 109617 274923
rect 107475 272117 108063 272151
rect 106997 272009 107175 272043
rect 106935 271819 106969 271959
rect 107203 271819 107237 271959
rect 106997 271735 107175 271769
rect 107413 271747 107447 272067
rect 108091 271747 108125 272067
rect 107475 271663 108063 271697
rect 107185 271501 108361 271535
rect 107101 271327 107135 271473
rect 108411 271327 108445 271473
rect 107185 271265 108361 271299
rect 107185 271131 108361 271165
rect 107101 270957 107135 271103
rect 108411 270957 108445 271103
rect 107185 270895 108361 270929
rect 108976 270837 109077 271005
rect 109456 272473 109494 272507
rect 109394 270718 109428 272414
rect 109522 270718 109556 272414
rect 109456 270625 109494 270659
rect 111536 280832 112612 280866
rect 111452 280676 111486 280804
rect 112662 280676 112696 280804
rect 111536 280614 112612 280648
rect 112982 280840 114058 280874
rect 112898 280644 112932 280812
rect 114108 280644 114142 280812
rect 112982 280582 114058 280616
rect 111536 280472 112612 280506
rect 111452 280316 111486 280444
rect 112662 280316 112696 280444
rect 111536 280254 112612 280288
rect 112982 280416 114058 280450
rect 112898 280220 112932 280388
rect 114108 280220 114142 280388
rect 112982 280158 114058 280192
rect 111536 280112 112612 280146
rect 111452 279956 111486 280084
rect 112662 279956 112696 280084
rect 111536 279894 112612 279928
rect 113012 280014 114088 280048
rect 112928 279938 112962 279986
rect 114138 279938 114172 279986
rect 113012 279876 114088 279910
rect 114342 279893 114377 279976
rect 111536 279752 112612 279786
rect 111452 279596 111486 279724
rect 112662 279596 112696 279724
rect 113012 279716 114088 279750
rect 112928 279640 112962 279688
rect 114138 279640 114172 279688
rect 113012 279578 114088 279612
rect 111536 279534 112612 279568
rect 114010 279348 114237 279417
rect 114669 280815 114845 280849
rect 114576 280419 114610 280787
rect 114904 280419 114938 280787
rect 114669 280357 114845 280391
rect 114885 280226 114948 280294
rect 114669 280129 114845 280163
rect 114576 279973 114610 280101
rect 114904 279973 114938 280101
rect 114669 279911 114845 279945
rect 114868 279813 114965 279861
rect 114669 279721 114845 279755
rect 114576 279565 114610 279693
rect 114904 279565 114938 279693
rect 114669 279503 114845 279537
rect 115360 280815 115536 280849
rect 115267 280419 115301 280787
rect 115595 280419 115629 280787
rect 115360 280357 115536 280391
rect 115257 280226 115320 280294
rect 115360 280129 115536 280163
rect 115267 279973 115301 280101
rect 115595 279973 115629 280101
rect 115360 279911 115536 279945
rect 115240 279813 115337 279861
rect 115360 279721 115536 279755
rect 115267 279565 115301 279693
rect 115595 279565 115629 279693
rect 115360 279503 115536 279537
rect 116147 280840 117223 280874
rect 116063 280644 116097 280812
rect 117273 280644 117307 280812
rect 116147 280582 117223 280616
rect 117593 280832 118669 280866
rect 117509 280676 117543 280804
rect 118719 280676 118753 280804
rect 117593 280614 118669 280648
rect 116147 280416 117223 280450
rect 116063 280220 116097 280388
rect 117273 280220 117307 280388
rect 116147 280158 117223 280192
rect 117593 280472 118669 280506
rect 117509 280316 117543 280444
rect 118719 280316 118753 280444
rect 117593 280254 118669 280288
rect 116117 280014 117193 280048
rect 115828 279893 115863 279976
rect 116033 279938 116067 279986
rect 117243 279938 117277 279986
rect 116117 279876 117193 279910
rect 117593 280112 118669 280146
rect 117509 279956 117543 280084
rect 118719 279956 118753 280084
rect 117593 279894 118669 279928
rect 117593 279752 118669 279786
rect 116117 279716 117193 279750
rect 116033 279640 116067 279688
rect 117243 279640 117277 279688
rect 116117 279578 117193 279612
rect 117509 279596 117543 279724
rect 118719 279596 118753 279724
rect 117593 279534 118669 279568
rect 115968 279348 116195 279417
rect 111536 279166 112612 279200
rect 111452 279010 111486 279138
rect 112662 279010 112696 279138
rect 111536 278948 112612 278982
rect 112982 279174 114058 279208
rect 112898 278978 112932 279146
rect 114108 278978 114142 279146
rect 112982 278916 114058 278950
rect 111536 278806 112612 278840
rect 111452 278650 111486 278778
rect 112662 278650 112696 278778
rect 111536 278588 112612 278622
rect 112982 278750 114058 278784
rect 112898 278554 112932 278722
rect 114108 278554 114142 278722
rect 112982 278492 114058 278526
rect 111536 278446 112612 278480
rect 111452 278290 111486 278418
rect 112662 278290 112696 278418
rect 111536 278228 112612 278262
rect 113012 278348 114088 278382
rect 112928 278272 112962 278320
rect 114138 278272 114172 278320
rect 113012 278210 114088 278244
rect 114342 278227 114377 278310
rect 111536 278086 112612 278120
rect 111452 277930 111486 278058
rect 112662 277930 112696 278058
rect 113012 278050 114088 278084
rect 112928 277974 112962 278022
rect 114138 277974 114172 278022
rect 113012 277912 114088 277946
rect 111536 277868 112612 277902
rect 114010 277682 114237 277751
rect 114669 279149 114845 279183
rect 114576 278753 114610 279121
rect 114904 278753 114938 279121
rect 114669 278691 114845 278725
rect 114885 278560 114948 278628
rect 114669 278463 114845 278497
rect 114576 278307 114610 278435
rect 114904 278307 114938 278435
rect 114669 278245 114845 278279
rect 114868 278147 114965 278195
rect 114669 278055 114845 278089
rect 114576 277899 114610 278027
rect 114904 277899 114938 278027
rect 114669 277837 114845 277871
rect 115360 279149 115536 279183
rect 115267 278753 115301 279121
rect 115595 278753 115629 279121
rect 115360 278691 115536 278725
rect 115257 278560 115320 278628
rect 115360 278463 115536 278497
rect 115267 278307 115301 278435
rect 115595 278307 115629 278435
rect 115360 278245 115536 278279
rect 115240 278147 115337 278195
rect 115360 278055 115536 278089
rect 115267 277899 115301 278027
rect 115595 277899 115629 278027
rect 115360 277837 115536 277871
rect 116147 279174 117223 279208
rect 116063 278978 116097 279146
rect 117273 278978 117307 279146
rect 116147 278916 117223 278950
rect 117593 279166 118669 279200
rect 117509 279010 117543 279138
rect 118719 279010 118753 279138
rect 117593 278948 118669 278982
rect 116147 278750 117223 278784
rect 116063 278554 116097 278722
rect 117273 278554 117307 278722
rect 116147 278492 117223 278526
rect 117593 278806 118669 278840
rect 117509 278650 117543 278778
rect 118719 278650 118753 278778
rect 117593 278588 118669 278622
rect 116117 278348 117193 278382
rect 115828 278227 115863 278310
rect 116033 278272 116067 278320
rect 117243 278272 117277 278320
rect 116117 278210 117193 278244
rect 117593 278446 118669 278480
rect 117509 278290 117543 278418
rect 118719 278290 118753 278418
rect 117593 278228 118669 278262
rect 117593 278086 118669 278120
rect 116117 278050 117193 278084
rect 116033 277974 116067 278022
rect 117243 277974 117277 278022
rect 116117 277912 117193 277946
rect 117509 277930 117543 278058
rect 118719 277930 118753 278058
rect 117593 277868 118669 277902
rect 115968 277682 116195 277751
rect 111536 277500 112612 277534
rect 111452 277344 111486 277472
rect 112662 277344 112696 277472
rect 111536 277282 112612 277316
rect 112982 277508 114058 277542
rect 112898 277312 112932 277480
rect 114108 277312 114142 277480
rect 112982 277250 114058 277284
rect 111536 277140 112612 277174
rect 111452 276984 111486 277112
rect 112662 276984 112696 277112
rect 111536 276922 112612 276956
rect 112982 277084 114058 277118
rect 112898 276888 112932 277056
rect 114108 276888 114142 277056
rect 112982 276826 114058 276860
rect 111536 276780 112612 276814
rect 111452 276624 111486 276752
rect 112662 276624 112696 276752
rect 111536 276562 112612 276596
rect 113012 276682 114088 276716
rect 112928 276606 112962 276654
rect 114138 276606 114172 276654
rect 113012 276544 114088 276578
rect 114342 276561 114377 276644
rect 111536 276420 112612 276454
rect 111452 276264 111486 276392
rect 112662 276264 112696 276392
rect 113012 276384 114088 276418
rect 112928 276308 112962 276356
rect 114138 276308 114172 276356
rect 113012 276246 114088 276280
rect 111536 276202 112612 276236
rect 114010 276016 114237 276085
rect 114669 277483 114845 277517
rect 114576 277087 114610 277455
rect 114904 277087 114938 277455
rect 114669 277025 114845 277059
rect 114885 276894 114948 276962
rect 114669 276797 114845 276831
rect 114576 276641 114610 276769
rect 114904 276641 114938 276769
rect 114669 276579 114845 276613
rect 114868 276481 114965 276529
rect 114669 276389 114845 276423
rect 114576 276233 114610 276361
rect 114904 276233 114938 276361
rect 114669 276171 114845 276205
rect 115360 277483 115536 277517
rect 115267 277087 115301 277455
rect 115595 277087 115629 277455
rect 115360 277025 115536 277059
rect 115257 276894 115320 276962
rect 115360 276797 115536 276831
rect 115267 276641 115301 276769
rect 115595 276641 115629 276769
rect 115360 276579 115536 276613
rect 115240 276481 115337 276529
rect 115360 276389 115536 276423
rect 115267 276233 115301 276361
rect 115595 276233 115629 276361
rect 115360 276171 115536 276205
rect 116147 277508 117223 277542
rect 116063 277312 116097 277480
rect 117273 277312 117307 277480
rect 116147 277250 117223 277284
rect 117593 277500 118669 277534
rect 117509 277344 117543 277472
rect 118719 277344 118753 277472
rect 117593 277282 118669 277316
rect 116147 277084 117223 277118
rect 116063 276888 116097 277056
rect 117273 276888 117307 277056
rect 116147 276826 117223 276860
rect 117593 277140 118669 277174
rect 117509 276984 117543 277112
rect 118719 276984 118753 277112
rect 117593 276922 118669 276956
rect 116117 276682 117193 276716
rect 115828 276561 115863 276644
rect 116033 276606 116067 276654
rect 117243 276606 117277 276654
rect 116117 276544 117193 276578
rect 117593 276780 118669 276814
rect 117509 276624 117543 276752
rect 118719 276624 118753 276752
rect 117593 276562 118669 276596
rect 117593 276420 118669 276454
rect 116117 276384 117193 276418
rect 116033 276308 116067 276356
rect 117243 276308 117277 276356
rect 116117 276246 117193 276280
rect 117509 276264 117543 276392
rect 118719 276264 118753 276392
rect 117593 276202 118669 276236
rect 115968 276016 116195 276085
rect 111536 275834 112612 275868
rect 111452 275678 111486 275806
rect 112662 275678 112696 275806
rect 111536 275616 112612 275650
rect 112982 275842 114058 275876
rect 112898 275646 112932 275814
rect 114108 275646 114142 275814
rect 112982 275584 114058 275618
rect 111536 275474 112612 275508
rect 111452 275318 111486 275446
rect 112662 275318 112696 275446
rect 111536 275256 112612 275290
rect 112982 275418 114058 275452
rect 112898 275222 112932 275390
rect 114108 275222 114142 275390
rect 112982 275160 114058 275194
rect 111536 275114 112612 275148
rect 111452 274958 111486 275086
rect 112662 274958 112696 275086
rect 111536 274896 112612 274930
rect 113012 275016 114088 275050
rect 112928 274940 112962 274988
rect 114138 274940 114172 274988
rect 113012 274878 114088 274912
rect 114342 274895 114377 274978
rect 111536 274754 112612 274788
rect 111452 274598 111486 274726
rect 112662 274598 112696 274726
rect 113012 274718 114088 274752
rect 112928 274642 112962 274690
rect 114138 274642 114172 274690
rect 113012 274580 114088 274614
rect 111536 274536 112612 274570
rect 114010 274350 114237 274419
rect 114669 275817 114845 275851
rect 114576 275421 114610 275789
rect 114904 275421 114938 275789
rect 114669 275359 114845 275393
rect 114885 275228 114948 275296
rect 114669 275131 114845 275165
rect 114576 274975 114610 275103
rect 114904 274975 114938 275103
rect 114669 274913 114845 274947
rect 114868 274815 114965 274863
rect 114669 274723 114845 274757
rect 114576 274567 114610 274695
rect 114904 274567 114938 274695
rect 114669 274505 114845 274539
rect 115360 275817 115536 275851
rect 115267 275421 115301 275789
rect 115595 275421 115629 275789
rect 115360 275359 115536 275393
rect 115257 275228 115320 275296
rect 115360 275131 115536 275165
rect 115267 274975 115301 275103
rect 115595 274975 115629 275103
rect 115360 274913 115536 274947
rect 115240 274815 115337 274863
rect 115360 274723 115536 274757
rect 115267 274567 115301 274695
rect 115595 274567 115629 274695
rect 115360 274505 115536 274539
rect 116147 275842 117223 275876
rect 116063 275646 116097 275814
rect 117273 275646 117307 275814
rect 116147 275584 117223 275618
rect 117593 275834 118669 275868
rect 117509 275678 117543 275806
rect 118719 275678 118753 275806
rect 117593 275616 118669 275650
rect 116147 275418 117223 275452
rect 116063 275222 116097 275390
rect 117273 275222 117307 275390
rect 116147 275160 117223 275194
rect 117593 275474 118669 275508
rect 117509 275318 117543 275446
rect 118719 275318 118753 275446
rect 117593 275256 118669 275290
rect 116117 275016 117193 275050
rect 115828 274895 115863 274978
rect 116033 274940 116067 274988
rect 117243 274940 117277 274988
rect 116117 274878 117193 274912
rect 117593 275114 118669 275148
rect 117509 274958 117543 275086
rect 118719 274958 118753 275086
rect 117593 274896 118669 274930
rect 117593 274754 118669 274788
rect 116117 274718 117193 274752
rect 116033 274642 116067 274690
rect 117243 274642 117277 274690
rect 116117 274580 117193 274614
rect 117509 274598 117543 274726
rect 118719 274598 118753 274726
rect 117593 274536 118669 274570
rect 115968 274350 116195 274419
rect 111536 274168 112612 274202
rect 111452 274012 111486 274140
rect 112662 274012 112696 274140
rect 111536 273950 112612 273984
rect 112982 274176 114058 274210
rect 112898 273980 112932 274148
rect 114108 273980 114142 274148
rect 112982 273918 114058 273952
rect 111536 273808 112612 273842
rect 111452 273652 111486 273780
rect 112662 273652 112696 273780
rect 111536 273590 112612 273624
rect 112982 273752 114058 273786
rect 112898 273556 112932 273724
rect 114108 273556 114142 273724
rect 112982 273494 114058 273528
rect 111536 273448 112612 273482
rect 111452 273292 111486 273420
rect 112662 273292 112696 273420
rect 111536 273230 112612 273264
rect 113012 273350 114088 273384
rect 112928 273274 112962 273322
rect 114138 273274 114172 273322
rect 113012 273212 114088 273246
rect 114342 273229 114377 273312
rect 111536 273088 112612 273122
rect 111452 272932 111486 273060
rect 112662 272932 112696 273060
rect 113012 273052 114088 273086
rect 112928 272976 112962 273024
rect 114138 272976 114172 273024
rect 113012 272914 114088 272948
rect 111536 272870 112612 272904
rect 114010 272684 114237 272753
rect 114669 274151 114845 274185
rect 114576 273755 114610 274123
rect 114904 273755 114938 274123
rect 114669 273693 114845 273727
rect 114885 273562 114948 273630
rect 114669 273465 114845 273499
rect 114576 273309 114610 273437
rect 114904 273309 114938 273437
rect 114669 273247 114845 273281
rect 114868 273149 114965 273197
rect 114669 273057 114845 273091
rect 114576 272901 114610 273029
rect 114904 272901 114938 273029
rect 114669 272839 114845 272873
rect 115360 274151 115536 274185
rect 115267 273755 115301 274123
rect 115595 273755 115629 274123
rect 115360 273693 115536 273727
rect 115257 273562 115320 273630
rect 115360 273465 115536 273499
rect 115267 273309 115301 273437
rect 115595 273309 115629 273437
rect 115360 273247 115536 273281
rect 115240 273149 115337 273197
rect 115360 273057 115536 273091
rect 115267 272901 115301 273029
rect 115595 272901 115629 273029
rect 115360 272839 115536 272873
rect 114982 272765 115027 272793
rect 115027 272765 115061 272793
rect 115061 272765 115144 272793
rect 115144 272765 115178 272793
rect 115178 272765 115228 272793
rect 114982 272739 115228 272765
rect 116147 274176 117223 274210
rect 116063 273980 116097 274148
rect 117273 273980 117307 274148
rect 116147 273918 117223 273952
rect 117593 274168 118669 274202
rect 117509 274012 117543 274140
rect 118719 274012 118753 274140
rect 117593 273950 118669 273984
rect 116147 273752 117223 273786
rect 116063 273556 116097 273724
rect 117273 273556 117307 273724
rect 116147 273494 117223 273528
rect 117593 273808 118669 273842
rect 117509 273652 117543 273780
rect 118719 273652 118753 273780
rect 117593 273590 118669 273624
rect 116117 273350 117193 273384
rect 115828 273229 115863 273312
rect 116033 273274 116067 273322
rect 117243 273274 117277 273322
rect 116117 273212 117193 273246
rect 117593 273448 118669 273482
rect 117509 273292 117543 273420
rect 118719 273292 118753 273420
rect 117593 273230 118669 273264
rect 117593 273088 118669 273122
rect 116117 273052 117193 273086
rect 116033 272976 116067 273024
rect 117243 272976 117277 273024
rect 116117 272914 117193 272948
rect 117509 272932 117543 273060
rect 118719 272932 118753 273060
rect 117593 272870 118669 272904
rect 114982 272705 115001 272739
rect 115001 272705 115204 272739
rect 115204 272705 115228 272739
rect 114982 272417 115228 272705
rect 115968 272684 116195 272753
rect 116628 272127 118134 272226
rect 113840 271699 114065 272014
rect 115017 271918 115559 272016
rect 113091 271540 113431 271629
rect 112594 271353 112722 271387
rect 112994 271353 113122 271387
rect 113394 271353 113522 271387
rect 113794 271353 113922 271387
rect 112532 271118 112566 271294
rect 112750 271118 112784 271294
rect 112932 271118 112966 271294
rect 113150 271118 113184 271294
rect 113332 271118 113366 271294
rect 113550 271118 113584 271294
rect 113732 271118 113766 271294
rect 113950 271118 113984 271294
rect 112594 271025 112722 271059
rect 112994 271025 113122 271059
rect 113394 271025 113522 271059
rect 113794 271025 113922 271059
rect 114653 271324 114781 271358
rect 114591 271089 114625 271265
rect 115053 271324 115181 271358
rect 114809 271089 114843 271265
rect 114991 271089 115025 271265
rect 115209 271089 115243 271265
rect 114653 270996 114781 271030
rect 115053 270996 115181 271030
rect 115897 271962 116025 271996
rect 116297 271962 116425 271996
rect 116697 271962 116825 271996
rect 117097 271962 117225 271996
rect 117497 271962 117625 271996
rect 117897 271962 118025 271996
rect 118297 271962 118425 271996
rect 118697 271962 118825 271996
rect 115835 270836 115869 271912
rect 116053 270836 116087 271912
rect 116235 270836 116269 271912
rect 116453 270836 116487 271912
rect 116635 270836 116669 271912
rect 116853 270836 116887 271912
rect 117035 270836 117069 271912
rect 117253 270836 117287 271912
rect 117435 270836 117469 271912
rect 117653 270836 117687 271912
rect 117835 270836 117869 271912
rect 118053 270836 118087 271912
rect 118235 270836 118269 271912
rect 118453 270836 118487 271912
rect 118635 270836 118669 271912
rect 118853 270836 118887 271912
rect 115897 270752 116025 270786
rect 116297 270752 116425 270786
rect 116697 270752 116825 270786
rect 117097 270752 117225 270786
rect 117497 270752 117625 270786
rect 117897 270752 118025 270786
rect 118297 270752 118425 270786
rect 118697 270752 118825 270786
rect 114086 270576 114501 270673
rect 112576 270262 112704 270296
rect 112976 270262 113104 270296
rect 113376 270262 113504 270296
rect 113776 270262 113904 270296
rect 114176 270262 114304 270296
rect 114576 270262 114704 270296
rect 114976 270262 115104 270296
rect 115376 270262 115504 270296
rect 115776 270262 115904 270296
rect 116176 270262 116304 270296
rect 116576 270262 116704 270296
rect 116976 270262 117104 270296
rect 117376 270262 117504 270296
rect 117776 270262 117904 270296
rect 118176 270262 118304 270296
rect 118576 270262 118704 270296
rect 112514 269136 112548 270212
rect 112732 269136 112766 270212
rect 112914 269136 112948 270212
rect 113132 269136 113166 270212
rect 113314 269136 113348 270212
rect 113532 269136 113566 270212
rect 113714 269136 113748 270212
rect 113932 269136 113966 270212
rect 114114 269136 114148 270212
rect 114332 269136 114366 270212
rect 114514 269136 114548 270212
rect 114732 269136 114766 270212
rect 114914 269136 114948 270212
rect 115132 269136 115166 270212
rect 115314 269136 115348 270212
rect 115532 269136 115566 270212
rect 115714 269136 115748 270212
rect 115932 269136 115966 270212
rect 116114 269136 116148 270212
rect 116332 269136 116366 270212
rect 116514 269136 116548 270212
rect 116732 269136 116766 270212
rect 116914 269136 116948 270212
rect 117132 269136 117166 270212
rect 117314 269136 117348 270212
rect 117532 269136 117566 270212
rect 117714 269136 117748 270212
rect 117932 269136 117966 270212
rect 118114 269136 118148 270212
rect 118332 269136 118366 270212
rect 118514 269136 118548 270212
rect 118732 269136 118766 270212
rect 112576 269052 112704 269086
rect 112976 269052 113104 269086
rect 113376 269052 113504 269086
rect 113776 269052 113904 269086
rect 114176 269052 114304 269086
rect 114576 269052 114704 269086
rect 114976 269052 115104 269086
rect 115376 269052 115504 269086
rect 115776 269052 115904 269086
rect 116176 269052 116304 269086
rect 116576 269052 116704 269086
rect 116976 269052 117104 269086
rect 117376 269052 117504 269086
rect 117776 269052 117904 269086
rect 118176 269052 118304 269086
rect 118576 269052 118704 269086
rect 114322 268826 117498 268883
rect 114322 268747 117498 268826
rect 120445 280684 120813 280718
rect 120383 280549 120417 280625
rect 120841 280549 120875 280625
rect 121145 280684 121513 280718
rect 121083 280549 121117 280625
rect 121541 280549 121575 280625
rect 120445 280456 120813 280490
rect 121145 280456 121513 280490
rect 120445 280300 120813 280334
rect 121145 280300 121513 280334
rect 120383 279765 120417 280241
rect 120841 279765 120875 280241
rect 121083 279765 121117 280241
rect 121541 279765 121575 280241
rect 120445 279672 120813 279706
rect 121145 279672 121513 279706
rect 120445 279516 120813 279550
rect 121145 279516 121513 279550
rect 120383 278981 120417 279457
rect 120841 278981 120875 279457
rect 121083 278981 121117 279457
rect 121541 278981 121575 279457
rect 120445 278888 120813 278922
rect 121145 278888 121513 278922
rect 120445 278732 120813 278766
rect 121145 278732 121513 278766
rect 120383 278197 120417 278673
rect 120841 278197 120875 278673
rect 121083 278197 121117 278673
rect 121541 278197 121575 278673
rect 120445 278104 120813 278138
rect 121145 278104 121513 278138
rect 120445 277948 120813 277982
rect 121145 277948 121513 277982
rect 120383 277413 120417 277889
rect 120841 277413 120875 277889
rect 121083 277413 121117 277889
rect 121541 277413 121575 277889
rect 120445 277320 120813 277354
rect 121145 277320 121513 277354
rect 120445 277164 120813 277198
rect 121145 277164 121513 277198
rect 120383 276629 120417 277105
rect 120841 276629 120875 277105
rect 121083 276629 121117 277105
rect 121541 276629 121575 277105
rect 120445 276536 120813 276570
rect 121145 276536 121513 276570
rect 120445 276380 120813 276414
rect 121145 276380 121513 276414
rect 120383 275845 120417 276321
rect 120841 275845 120875 276321
rect 120958 276054 121014 276118
rect 121083 275845 121117 276321
rect 121541 275845 121575 276321
rect 120445 275752 120813 275786
rect 121145 275752 121513 275786
rect 120445 275596 120813 275630
rect 121145 275596 121513 275630
rect 120383 275061 120417 275537
rect 120841 275061 120875 275537
rect 120445 274968 120813 275002
rect 120445 274812 120813 274846
rect 120383 274277 120417 274753
rect 120841 274277 120875 274753
rect 121083 275061 121117 275537
rect 121541 275061 121575 275537
rect 121145 274968 121513 275002
rect 121145 274812 121513 274846
rect 121083 274277 121117 274753
rect 121541 274277 121575 274753
rect 120445 274184 120813 274218
rect 121145 274184 121513 274218
rect 120445 274028 120813 274062
rect 121145 274028 121513 274062
rect 120383 273493 120417 273969
rect 120841 273493 120875 273969
rect 120961 273692 121017 273756
rect 121083 273493 121117 273969
rect 121541 273493 121575 273969
rect 120445 273400 120813 273434
rect 121145 273400 121513 273434
rect 120445 273244 120813 273278
rect 121145 273244 121513 273278
rect 120383 272709 120417 273185
rect 120841 272709 120875 273185
rect 121083 272709 121117 273185
rect 121541 272709 121575 273185
rect 120445 272616 120813 272650
rect 121145 272616 121513 272650
rect 120445 272460 120813 272494
rect 121145 272460 121513 272494
rect 120383 271925 120417 272401
rect 120841 271925 120875 272401
rect 121083 271925 121117 272401
rect 121541 271925 121575 272401
rect 120445 271832 120813 271866
rect 121145 271832 121513 271866
rect 120445 271676 120813 271710
rect 121145 271676 121513 271710
rect 120383 271141 120417 271617
rect 120841 271141 120875 271617
rect 121083 271141 121117 271617
rect 121541 271141 121575 271617
rect 120445 271048 120813 271082
rect 121145 271048 121513 271082
rect 120445 270892 120813 270926
rect 121145 270892 121513 270926
rect 120383 270357 120417 270833
rect 120841 270357 120875 270833
rect 121083 270357 121117 270833
rect 121541 270357 121575 270833
rect 120445 270264 120813 270298
rect 121145 270264 121513 270298
rect 120445 270108 120813 270142
rect 121145 270108 121513 270142
rect 120383 269573 120417 270049
rect 120841 269573 120875 270049
rect 121083 269573 121117 270049
rect 121541 269573 121575 270049
rect 120445 269480 120813 269514
rect 121145 269480 121513 269514
rect 120445 269324 120813 269358
rect 121145 269324 121513 269358
rect 120383 269189 120417 269265
rect 120841 269189 120875 269265
rect 120445 269096 120813 269130
rect 121083 269189 121117 269265
rect 121541 269189 121575 269265
rect 121145 269096 121513 269130
rect 122372 280470 122740 280504
rect 123072 280470 123440 280504
rect 122310 279935 122344 280411
rect 122768 279935 122802 280411
rect 123010 279935 123044 280411
rect 123468 279935 123502 280411
rect 121849 279275 122178 279887
rect 122178 279275 122191 279887
rect 122372 279842 122740 279876
rect 123072 279842 123440 279876
rect 122372 279686 122740 279720
rect 123072 279686 123440 279720
rect 122310 279151 122344 279627
rect 122768 279151 122802 279627
rect 123010 279151 123044 279627
rect 123468 279151 123502 279627
rect 122372 279058 122740 279092
rect 123072 279058 123440 279092
rect 122430 278313 123274 278347
rect 122368 277804 122402 278254
rect 123302 277804 123336 278254
rect 122430 277711 123274 277745
rect 122432 277547 123200 277581
rect 122370 277412 122404 277488
rect 123228 277412 123262 277488
rect 122432 277319 123200 277353
rect 123672 278127 124194 278161
rect 123610 277406 123644 278068
rect 124222 277406 124256 278068
rect 123672 277313 124194 277347
rect 123736 276881 123913 277034
rect 122454 276715 123816 276749
rect 122392 276504 122426 276656
rect 123844 276504 123878 276656
rect 122454 276411 123816 276445
rect 122120 276060 122144 276131
rect 122144 276060 122404 276131
rect 124465 275982 124549 276083
rect 122478 275823 122854 275857
rect 123114 275823 123490 275857
rect 123750 275823 124126 275857
rect 124386 275823 124762 275857
rect 122385 275727 122419 275795
rect 122913 275727 122947 275795
rect 123021 275727 123055 275795
rect 123549 275727 123583 275795
rect 123657 275727 123691 275795
rect 124185 275727 124219 275795
rect 124293 275727 124327 275795
rect 124821 275727 124855 275795
rect 122478 275665 122854 275699
rect 123114 275665 123490 275699
rect 123750 275665 124126 275699
rect 124386 275665 124762 275699
rect 123245 275173 123426 275386
rect 122968 274900 123936 274934
rect 122906 274674 122940 274850
rect 123964 274674 123998 274850
rect 122968 274590 123936 274624
rect 122293 274316 122461 274350
rect 122709 274316 122877 274350
rect 123527 274408 123647 274445
rect 123125 274316 123293 274350
rect 123541 274316 123709 274350
rect 123957 274316 124125 274350
rect 122231 273790 122265 274266
rect 122489 273790 122523 274266
rect 122647 273790 122681 274266
rect 122905 273790 122939 274266
rect 123063 273790 123097 274266
rect 123321 273790 123355 274266
rect 123479 273790 123513 274266
rect 123737 273790 123771 274266
rect 123895 273790 123929 274266
rect 124153 273790 124187 274266
rect 124373 274316 124541 274350
rect 124311 273790 124345 274266
rect 124569 273790 124603 274266
rect 122293 273706 122461 273740
rect 122709 273706 122877 273740
rect 123125 273706 123293 273740
rect 123541 273706 123709 273740
rect 123957 273706 124125 273740
rect 124373 273706 124541 273740
rect 122141 272860 122509 272894
rect 122079 272725 122113 272801
rect 122537 272725 122571 272801
rect 122141 272632 122509 272666
rect 122841 272860 123209 272894
rect 122779 272725 122813 272801
rect 123237 272725 123271 272801
rect 122841 272632 123209 272666
rect 122141 272476 122509 272510
rect 122841 272476 123209 272510
rect 123355 272446 123444 272626
rect 122079 271941 122113 272417
rect 122537 271941 122571 272417
rect 122654 272150 122710 272214
rect 122779 271941 122813 272417
rect 123237 271941 123271 272417
rect 122141 271848 122509 271882
rect 122841 271848 123209 271882
rect 122141 271692 122509 271726
rect 122841 271692 123209 271726
rect 122079 271157 122113 271633
rect 122537 271157 122571 271633
rect 122141 271064 122509 271098
rect 122141 270908 122509 270942
rect 122079 270373 122113 270849
rect 122537 270373 122571 270849
rect 122779 271157 122813 271633
rect 123237 271157 123271 271633
rect 122841 271064 123209 271098
rect 122841 270908 123209 270942
rect 122779 270373 122813 270849
rect 123237 270373 123271 270849
rect 122141 270280 122509 270314
rect 122841 270280 123209 270314
rect 122141 270124 122509 270158
rect 122841 270124 123209 270158
rect 122079 269589 122113 270065
rect 122537 269589 122571 270065
rect 122657 269788 122713 269852
rect 122779 269589 122813 270065
rect 123237 269589 123271 270065
rect 122141 269496 122509 269530
rect 122841 269496 123209 269530
rect 122141 269340 122509 269374
rect 122079 269205 122113 269281
rect 122537 269205 122571 269281
rect 122141 269112 122509 269146
rect 122841 269340 123209 269374
rect 122779 269205 122813 269281
rect 123237 269205 123271 269281
rect 122841 269112 123209 269146
rect 124204 272532 124680 272566
rect 124120 272336 124154 272504
rect 124730 272336 124764 272504
rect 124204 272274 124680 272308
rect 124204 272116 124680 272150
rect 124120 271920 124154 272088
rect 124730 271920 124764 272088
rect 124204 271858 124680 271892
rect 124204 271700 124680 271734
rect 124120 271504 124154 271672
rect 124730 271504 124764 271672
rect 124204 271442 124680 271476
rect 124204 271284 124680 271318
rect 124120 271088 124154 271256
rect 124730 271088 124764 271256
rect 124204 271026 124680 271060
rect 124204 270868 124680 270902
rect 124120 270672 124154 270840
rect 124730 270672 124764 270840
rect 124204 270610 124680 270644
rect 124204 270452 124680 270486
rect 124120 270256 124154 270424
rect 124730 270256 124764 270424
rect 124204 270194 124680 270228
rect 124204 270036 124680 270070
rect 124120 269840 124154 270008
rect 124730 269840 124764 270008
rect 124204 269778 124680 269812
rect 124204 269620 124680 269654
rect 124120 269424 124154 269592
rect 124730 269424 124764 269592
rect 124204 269362 124680 269396
rect 125790 268342 128055 275158
<< metal1 >>
rect 105796 283673 113672 283895
rect 105796 282423 106140 283673
rect 113415 282909 113672 283673
rect 113415 282423 125337 282909
rect 105796 282251 125337 282423
rect 102098 281654 103259 281810
rect 102098 280847 102248 281654
rect 103117 281274 103259 281654
rect 103117 281095 108300 281274
rect 103117 280847 103259 281095
rect 108146 281064 108300 281095
rect 108146 280949 108295 281064
rect 102098 280720 103259 280847
rect 106361 280885 106485 280891
rect 106361 280851 106373 280885
rect 106473 280851 106485 280885
rect 106361 280845 106485 280851
rect 106761 280885 109685 280949
rect 106761 280851 106773 280885
rect 106873 280879 107173 280885
rect 106873 280851 106885 280879
rect 106761 280845 106885 280851
rect 107161 280851 107173 280879
rect 107273 280879 107573 280885
rect 107273 280851 107285 280879
rect 107161 280845 107285 280851
rect 107561 280851 107573 280879
rect 107673 280879 107973 280885
rect 107673 280851 107685 280879
rect 107561 280845 107685 280851
rect 107961 280851 107973 280879
rect 108073 280879 108373 280885
rect 108073 280851 108085 280879
rect 107961 280845 108085 280851
rect 108196 280813 108255 280879
rect 108361 280851 108373 280879
rect 108473 280879 108773 280885
rect 108473 280851 108485 280879
rect 108361 280845 108485 280851
rect 108761 280851 108773 280879
rect 108873 280879 109173 280885
rect 108873 280851 108885 280879
rect 108761 280845 108885 280851
rect 109161 280851 109173 280879
rect 109273 280879 109573 280885
rect 109273 280851 109285 280879
rect 109161 280845 109285 280851
rect 109561 280851 109573 280879
rect 109673 280851 109685 280885
rect 109561 280845 109685 280851
rect 109961 280885 110085 280891
rect 109961 280851 109973 280885
rect 110073 280851 110085 280885
rect 109961 280845 110085 280851
rect 106305 280801 106351 280813
rect 106305 279805 106311 280801
rect 106345 279805 106351 280801
rect 106305 279793 106351 279805
rect 106495 280801 106541 280813
rect 106495 279805 106501 280801
rect 106535 279805 106541 280801
rect 106495 279793 106541 279805
rect 106705 280801 106751 280813
rect 106705 279805 106711 280801
rect 106745 279805 106751 280801
rect 106705 279793 106751 279805
rect 106895 280801 106996 280813
rect 106895 279805 106901 280801
rect 106935 279805 106996 280801
rect 106895 279793 106996 279805
rect 107105 280801 107151 280813
rect 107105 279805 107111 280801
rect 107145 279805 107151 280801
rect 107105 279793 107151 279805
rect 107295 280801 107396 280813
rect 107295 279805 107301 280801
rect 107335 279805 107396 280801
rect 107295 279793 107396 279805
rect 107505 280801 107551 280813
rect 107505 279805 107511 280801
rect 107545 279805 107551 280801
rect 107505 279793 107551 279805
rect 107695 280801 107796 280813
rect 107695 279805 107701 280801
rect 107735 279805 107796 280801
rect 107695 279793 107796 279805
rect 107905 280801 107951 280813
rect 107905 279805 107911 280801
rect 107945 279805 107951 280801
rect 107905 279793 107951 279805
rect 108095 280801 108351 280813
rect 108095 279805 108101 280801
rect 108135 279805 108311 280801
rect 108345 279805 108351 280801
rect 108095 279793 108351 279805
rect 108495 280801 108541 280813
rect 108495 279805 108501 280801
rect 108535 279805 108541 280801
rect 108495 279793 108541 279805
rect 108650 280801 108751 280813
rect 108650 279805 108711 280801
rect 108745 279805 108751 280801
rect 108650 279793 108751 279805
rect 108895 280801 108941 280813
rect 108895 279805 108901 280801
rect 108935 279805 108941 280801
rect 108895 279793 108941 279805
rect 109050 280801 109151 280813
rect 109050 279805 109111 280801
rect 109145 279805 109151 280801
rect 109050 279793 109151 279805
rect 109295 280801 109341 280813
rect 109295 279805 109301 280801
rect 109335 279805 109341 280801
rect 109295 279793 109341 279805
rect 109450 280801 109551 280813
rect 109450 279805 109511 280801
rect 109545 279805 109551 280801
rect 109450 279793 109551 279805
rect 109695 280801 109741 280813
rect 109695 279805 109701 280801
rect 109735 279805 109741 280801
rect 109695 279793 109741 279805
rect 109905 280801 109951 280813
rect 109905 279805 109911 280801
rect 109945 279805 109951 280801
rect 109905 279793 109951 279805
rect 110095 280801 110141 280813
rect 110095 279805 110101 280801
rect 110135 279805 110141 280801
rect 110095 279793 110141 279805
rect 106361 279755 106485 279761
rect 106361 279721 106373 279755
rect 106473 279721 106485 279755
rect 106361 279715 106485 279721
rect 106761 279755 106885 279761
rect 106761 279721 106773 279755
rect 106873 279721 106885 279755
rect 106761 279715 106885 279721
rect 106941 279401 106996 279793
rect 107161 279755 107285 279761
rect 107161 279721 107173 279755
rect 107273 279721 107285 279755
rect 107161 279715 107285 279721
rect 107341 279642 107396 279793
rect 107561 279755 107685 279761
rect 107561 279721 107573 279755
rect 107673 279721 107685 279755
rect 107561 279715 107685 279721
rect 107741 279642 107796 279793
rect 107961 279755 108085 279761
rect 107961 279721 107973 279755
rect 108073 279721 108085 279755
rect 107961 279715 108085 279721
rect 108361 279755 108485 279761
rect 108361 279721 108373 279755
rect 108473 279721 108485 279755
rect 108361 279715 108485 279721
rect 107341 279599 107796 279642
rect 107341 279512 107422 279599
rect 107721 279519 107796 279599
rect 108650 279641 108705 279793
rect 108761 279755 108885 279761
rect 108761 279721 108773 279755
rect 108873 279721 108885 279755
rect 108761 279715 108885 279721
rect 109050 279641 109105 279793
rect 109161 279755 109285 279761
rect 109161 279721 109173 279755
rect 109273 279721 109285 279755
rect 109161 279715 109285 279721
rect 108650 279599 109105 279641
rect 108650 279519 108732 279599
rect 107721 279512 108732 279519
rect 109031 279512 109105 279599
rect 107341 279471 109105 279512
rect 109450 279401 109505 279793
rect 109561 279755 109685 279761
rect 109561 279721 109573 279755
rect 109673 279721 109685 279755
rect 109561 279715 109685 279721
rect 109961 279755 110085 279761
rect 109961 279721 109973 279755
rect 110073 279721 110085 279755
rect 109961 279715 110085 279721
rect 106941 279348 109505 279401
rect 107340 279238 107584 279258
rect 107340 279130 107381 279238
rect 106148 279108 107381 279130
rect 107553 279108 107584 279238
rect 106148 279065 107584 279108
rect 106148 279063 107582 279065
rect 106148 278530 106235 279063
rect 106368 279057 107582 279063
rect 106368 279023 106380 279057
rect 107570 279023 107582 279057
rect 106368 279017 107582 279023
rect 106281 278995 106327 279007
rect 106281 278773 106287 278995
rect 106321 278773 106327 278995
rect 106281 278761 106327 278773
rect 107623 278995 107669 279007
rect 107623 278773 107629 278995
rect 107663 278773 107669 278995
rect 107623 278761 107669 278773
rect 106368 278745 107582 278751
rect 106368 278711 106380 278745
rect 107570 278711 107582 278745
rect 106368 278705 107582 278711
rect 106368 278638 107796 278705
rect 106148 278463 107582 278530
rect 106368 278457 107582 278463
rect 106368 278423 106380 278457
rect 107570 278423 107582 278457
rect 106368 278417 107582 278423
rect 106281 278395 106327 278407
rect 104099 278379 106210 278382
rect 106281 278379 106287 278395
rect 104099 278179 106287 278379
rect 104099 278177 106210 278179
rect 102098 276478 103259 276621
rect 102098 275681 102261 276478
rect 103092 276209 103259 276478
rect 104099 276209 104304 278177
rect 106281 278173 106287 278179
rect 106321 278173 106327 278395
rect 106281 278161 106327 278173
rect 107623 278395 107669 278407
rect 107623 278173 107629 278395
rect 107663 278173 107669 278395
rect 107623 278161 107669 278173
rect 106368 278145 107582 278151
rect 106368 278111 106380 278145
rect 107570 278111 107582 278145
rect 106368 278105 107582 278111
rect 107709 278105 107796 278638
rect 106368 278068 107796 278105
rect 106368 278038 106941 278068
rect 103092 276004 104304 276209
rect 104854 277825 106544 277826
rect 104854 277627 106760 277825
rect 106902 277789 106941 278038
rect 107098 278038 107796 278068
rect 107098 277799 107130 278038
rect 107098 277789 107553 277799
rect 106902 277751 107553 277789
rect 106902 277724 107015 277751
rect 106957 277627 107015 277724
rect 104854 277449 107015 277627
rect 107487 277449 107553 277751
rect 104854 277407 107553 277449
rect 104854 277397 106760 277407
rect 106957 277403 107553 277407
rect 103092 275681 103259 276004
rect 102098 275531 103259 275681
rect 102557 274145 104316 274146
rect 104854 274145 105283 277397
rect 106959 277216 107081 277403
rect 106491 277210 107525 277216
rect 106491 277176 106503 277210
rect 107513 277176 107525 277210
rect 106491 277170 107525 277176
rect 106404 277148 106450 277160
rect 106404 277106 106410 277148
rect 106444 277106 106450 277148
rect 106404 276855 106450 277106
rect 107566 277158 107612 277160
rect 107566 277148 107889 277158
rect 107566 277106 107572 277148
rect 107606 277125 107889 277148
rect 107606 277106 107782 277125
rect 107566 277102 107782 277106
rect 107566 277094 107612 277102
rect 106491 277078 107525 277084
rect 106491 277044 106503 277078
rect 107513 277044 107525 277078
rect 106491 277038 107525 277044
rect 107754 276855 107782 277102
rect 106404 276842 107782 276855
rect 107861 276842 107889 277125
rect 106404 276808 107889 276842
rect 106294 276290 106623 276403
rect 106294 275337 106375 276290
rect 106100 274853 106375 275337
rect 106549 274853 106623 276290
rect 107947 276127 108079 276165
rect 107947 276009 107978 276127
rect 108049 276009 108079 276127
rect 107947 275882 108079 276009
rect 109196 275969 109291 279348
rect 109517 279089 110059 279151
rect 109517 277895 109569 279089
rect 109781 279083 110059 279089
rect 109781 279049 109793 279083
rect 110047 279049 110059 279083
rect 109781 279043 110059 279049
rect 109725 278999 109771 279011
rect 109725 278903 109731 278999
rect 109659 278872 109731 278903
rect 109659 278009 109692 278872
rect 109659 277985 109731 278009
rect 109765 277985 109771 278999
rect 109659 277973 109771 277985
rect 110069 278999 110165 279011
rect 110069 277985 110075 278999
rect 110109 278060 110165 278999
rect 110109 277985 110256 278060
rect 110069 277973 110256 277985
rect 109781 277935 110059 277941
rect 109781 277901 109793 277935
rect 110047 277901 110059 277935
rect 109781 277895 110059 277901
rect 109517 277833 110059 277895
rect 109517 277341 109569 277833
rect 109781 277827 110059 277833
rect 109781 277793 109793 277827
rect 110047 277793 110059 277827
rect 109781 277787 110059 277793
rect 110115 277755 110256 277973
rect 109413 277299 109569 277341
rect 109413 276623 109452 277299
rect 109533 276639 109569 277299
rect 109659 277743 109771 277755
rect 109659 277718 109731 277743
rect 109659 276855 109687 277718
rect 109659 276825 109731 276855
rect 109725 276729 109731 276825
rect 109765 276729 109771 277743
rect 109725 276717 109771 276729
rect 110069 277743 110256 277755
rect 110069 276729 110075 277743
rect 110109 276729 110256 277743
rect 110069 276717 110256 276729
rect 109781 276679 110059 276685
rect 109781 276645 109793 276679
rect 110047 276645 110059 276679
rect 109781 276639 110059 276645
rect 109533 276623 110059 276639
rect 109413 276577 110059 276623
rect 110149 276420 110256 276717
rect 109824 276348 110271 276420
rect 109824 276166 109918 276348
rect 110180 276166 110271 276348
rect 109824 276093 110271 276166
rect 109193 275949 109712 275969
rect 107507 275832 109067 275882
rect 109193 275859 109262 275949
rect 109636 275859 109712 275949
rect 109193 275836 109712 275859
rect 107507 275765 107567 275832
rect 109007 275765 109067 275832
rect 106951 275759 107129 275765
rect 106951 275725 106963 275759
rect 107117 275725 107129 275759
rect 106951 275719 107129 275725
rect 107451 275759 107629 275765
rect 107451 275725 107463 275759
rect 107617 275725 107629 275759
rect 107451 275719 107629 275725
rect 107951 275759 108629 275765
rect 107951 275725 107963 275759
rect 108117 275727 108463 275759
rect 108117 275725 108227 275727
rect 107951 275719 108227 275725
rect 108129 275709 108227 275719
rect 106864 275697 106910 275709
rect 106864 274951 106870 275697
rect 106904 274951 106910 275697
rect 106864 274939 106910 274951
rect 107170 275697 107216 275709
rect 107170 274951 107176 275697
rect 107210 274951 107216 275697
rect 107170 274939 107216 274951
rect 107364 275697 107410 275709
rect 107364 274951 107370 275697
rect 107404 274951 107410 275697
rect 107364 274939 107410 274951
rect 107670 275697 107716 275709
rect 107670 274951 107676 275697
rect 107710 275393 107716 275697
rect 107864 275697 107910 275709
rect 107864 275393 107870 275697
rect 107710 275259 107870 275393
rect 107710 274951 107716 275259
rect 107670 274939 107716 274951
rect 107864 274951 107870 275259
rect 107904 274951 107910 275697
rect 107864 274939 107910 274951
rect 108170 275697 108227 275709
rect 108170 274951 108176 275697
rect 108210 275576 108227 275697
rect 108353 275725 108463 275727
rect 108617 275725 108629 275759
rect 108353 275719 108629 275725
rect 108951 275759 109129 275765
rect 108951 275725 108963 275759
rect 109117 275725 109129 275759
rect 108951 275719 109129 275725
rect 109451 275759 109629 275765
rect 109451 275725 109463 275759
rect 109617 275725 109629 275759
rect 109451 275719 109629 275725
rect 108353 275709 108451 275719
rect 108353 275697 108410 275709
rect 108353 275576 108370 275697
rect 108210 275522 108370 275576
rect 108210 275393 108216 275522
rect 108364 275393 108370 275522
rect 108210 275259 108370 275393
rect 108210 274951 108216 275259
rect 108170 274939 108216 274951
rect 108364 274951 108370 275259
rect 108404 274951 108410 275697
rect 108364 274939 108410 274951
rect 108670 275697 108716 275709
rect 108670 274951 108676 275697
rect 108710 275393 108716 275697
rect 108864 275697 108910 275709
rect 108864 275393 108870 275697
rect 108710 275259 108870 275393
rect 108710 274951 108716 275259
rect 108670 274939 108716 274951
rect 108864 274951 108870 275259
rect 108904 274951 108910 275697
rect 108864 274939 108910 274951
rect 109170 275697 109216 275709
rect 109170 274951 109176 275697
rect 109210 274951 109216 275697
rect 109170 274939 109216 274951
rect 109364 275697 109410 275709
rect 109364 274951 109370 275697
rect 109404 274951 109410 275697
rect 109364 274939 109410 274951
rect 109670 275697 109716 275709
rect 109670 274951 109676 275697
rect 109710 274951 109716 275697
rect 109670 274939 109716 274951
rect 106951 274923 107129 274929
rect 106951 274889 106963 274923
rect 107117 274889 107129 274923
rect 106951 274883 107129 274889
rect 107451 274923 107629 274929
rect 107451 274889 107463 274923
rect 107617 274889 107629 274923
rect 107451 274883 107629 274889
rect 107951 274923 108129 274929
rect 107951 274889 107963 274923
rect 108117 274889 108129 274923
rect 107951 274883 108129 274889
rect 108451 274923 108629 274929
rect 108451 274889 108463 274923
rect 108617 274889 108629 274923
rect 108451 274883 108629 274889
rect 108951 274923 109129 274929
rect 108951 274889 108963 274923
rect 109117 274889 109129 274923
rect 108951 274883 109129 274889
rect 109451 274923 109629 274929
rect 109451 274889 109463 274923
rect 109617 274889 109629 274923
rect 109451 274883 109629 274889
rect 106100 274731 106623 274853
rect 106100 274505 106622 274731
rect 110521 274509 111012 282251
rect 119259 281225 119845 282251
rect 119257 281145 119845 281225
rect 112970 280874 114070 280880
rect 111524 280866 112624 280872
rect 111524 280832 111536 280866
rect 112612 280832 112624 280866
rect 112970 280840 112982 280874
rect 114058 280840 114070 280874
rect 116135 280874 117235 280880
rect 112970 280834 114070 280840
rect 114657 280849 114857 280855
rect 111524 280826 112624 280832
rect 111404 280804 111492 280816
rect 111404 280676 111452 280804
rect 111486 280676 111492 280804
rect 111404 280664 111492 280676
rect 112656 280804 112744 280816
rect 112656 280676 112662 280804
rect 112696 280748 112744 280804
rect 112850 280812 112938 280824
rect 112850 280748 112898 280812
rect 112696 280686 112898 280748
rect 112696 280676 112744 280686
rect 112656 280664 112744 280676
rect 111404 280456 111446 280664
rect 111524 280648 112624 280654
rect 111524 280614 111536 280648
rect 112612 280614 112624 280648
rect 111524 280608 112624 280614
rect 112702 280632 112744 280664
rect 112850 280644 112898 280686
rect 112932 280644 112938 280812
rect 112850 280632 112938 280644
rect 114102 280812 114190 280824
rect 114102 280644 114108 280812
rect 114142 280758 114190 280812
rect 114657 280815 114669 280849
rect 114845 280815 114857 280849
rect 114657 280809 114857 280815
rect 115348 280849 115548 280855
rect 115348 280815 115360 280849
rect 115536 280815 115548 280849
rect 116135 280840 116147 280874
rect 117223 280840 117235 280874
rect 116135 280834 117235 280840
rect 117581 280866 118681 280872
rect 117581 280832 117593 280866
rect 118669 280832 118681 280866
rect 117581 280826 118681 280832
rect 115348 280809 115548 280815
rect 116015 280812 116103 280824
rect 114570 280787 114616 280799
rect 114570 280758 114576 280787
rect 114142 280644 114576 280758
rect 114102 280632 114576 280644
rect 111524 280506 112624 280512
rect 111524 280472 111536 280506
rect 112612 280472 112624 280506
rect 111524 280466 112624 280472
rect 112702 280456 112746 280632
rect 111404 280444 111492 280456
rect 111404 280316 111452 280444
rect 111486 280316 111492 280444
rect 111404 280304 111492 280316
rect 112656 280444 112746 280456
rect 112656 280316 112662 280444
rect 112696 280412 112746 280444
rect 112850 280532 112892 280632
rect 114148 280625 114576 280632
rect 112970 280616 114070 280622
rect 112970 280582 112982 280616
rect 114058 280582 114070 280616
rect 112970 280576 114070 280582
rect 114148 280532 114190 280625
rect 112850 280494 114190 280532
rect 112696 280364 112744 280412
rect 112850 280400 112892 280494
rect 112970 280450 114070 280456
rect 112970 280416 112982 280450
rect 114058 280416 114070 280450
rect 112970 280410 114070 280416
rect 114148 280400 114190 280494
rect 114570 280419 114576 280625
rect 114610 280419 114616 280787
rect 114570 280407 114616 280419
rect 114898 280787 114944 280799
rect 114898 280419 114904 280787
rect 114938 280419 114944 280787
rect 114898 280407 114944 280419
rect 115261 280787 115307 280799
rect 115261 280419 115267 280787
rect 115301 280419 115307 280787
rect 115261 280407 115307 280419
rect 115589 280787 115635 280799
rect 115589 280419 115595 280787
rect 115629 280758 115635 280787
rect 116015 280758 116063 280812
rect 115629 280644 116063 280758
rect 116097 280644 116103 280812
rect 115629 280632 116103 280644
rect 117267 280812 117355 280824
rect 117267 280644 117273 280812
rect 117307 280748 117355 280812
rect 117461 280804 117549 280816
rect 117461 280748 117509 280804
rect 117307 280686 117509 280748
rect 117307 280644 117355 280686
rect 117267 280632 117355 280644
rect 117461 280676 117509 280686
rect 117543 280676 117549 280804
rect 117461 280664 117549 280676
rect 118713 280804 118801 280816
rect 118713 280676 118719 280804
rect 118753 280676 118801 280804
rect 118713 280664 118801 280676
rect 117461 280632 117503 280664
rect 115629 280625 116057 280632
rect 115629 280419 115635 280625
rect 115589 280407 115635 280419
rect 116015 280532 116057 280625
rect 116135 280616 117235 280622
rect 116135 280582 116147 280616
rect 117223 280582 117235 280616
rect 116135 280576 117235 280582
rect 117313 280532 117355 280632
rect 116015 280494 117355 280532
rect 112850 280388 112938 280400
rect 112850 280364 112898 280388
rect 112696 280316 112898 280364
rect 112656 280304 112898 280316
rect 111404 280096 111446 280304
rect 112702 280302 112898 280304
rect 111524 280288 112624 280294
rect 111524 280254 111536 280288
rect 112612 280254 112624 280288
rect 111524 280248 112624 280254
rect 111524 280146 112624 280152
rect 111524 280112 111536 280146
rect 112612 280112 112624 280146
rect 111524 280106 112624 280112
rect 112702 280096 112744 280302
rect 112850 280220 112898 280302
rect 112932 280220 112938 280388
rect 112850 280208 112938 280220
rect 114102 280388 114190 280400
rect 116015 280400 116057 280494
rect 116135 280450 117235 280456
rect 116135 280416 116147 280450
rect 117223 280416 117235 280450
rect 116135 280410 117235 280416
rect 117313 280400 117355 280494
rect 117459 280456 117503 280632
rect 117581 280648 118681 280654
rect 117581 280614 117593 280648
rect 118669 280614 118681 280648
rect 117581 280608 118681 280614
rect 117581 280506 118681 280512
rect 117581 280472 117593 280506
rect 118669 280472 118681 280506
rect 117581 280466 118681 280472
rect 118759 280456 118801 280664
rect 117459 280444 117549 280456
rect 117459 280412 117509 280444
rect 114102 280220 114108 280388
rect 114142 280220 114190 280388
rect 114657 280391 114857 280397
rect 114657 280357 114669 280391
rect 114845 280357 114857 280391
rect 114657 280351 114857 280357
rect 115348 280391 115548 280397
rect 115348 280357 115360 280391
rect 115536 280357 115548 280391
rect 115348 280351 115548 280357
rect 116015 280388 116103 280400
rect 114720 280283 114790 280351
rect 114102 280208 114190 280220
rect 114308 280199 114790 280283
rect 114865 280294 114970 280311
rect 114865 280226 114885 280294
rect 114948 280226 114970 280294
rect 114865 280204 114970 280226
rect 115235 280294 115340 280311
rect 115235 280226 115257 280294
rect 115320 280226 115340 280294
rect 115235 280204 115340 280226
rect 115415 280283 115485 280351
rect 112970 280192 114070 280198
rect 112970 280158 112982 280192
rect 114058 280158 114070 280192
rect 112970 280152 114070 280158
rect 111404 280084 111492 280096
rect 111404 279956 111452 280084
rect 111486 279956 111492 280084
rect 111404 279944 111492 279956
rect 112656 280084 112744 280096
rect 114308 280084 114343 280199
rect 114720 280169 114790 280199
rect 115415 280199 115897 280283
rect 116015 280220 116063 280388
rect 116097 280220 116103 280388
rect 116015 280208 116103 280220
rect 117267 280388 117355 280400
rect 117267 280220 117273 280388
rect 117307 280364 117355 280388
rect 117461 280364 117509 280412
rect 117307 280316 117509 280364
rect 117543 280316 117549 280444
rect 117307 280304 117549 280316
rect 118713 280444 118801 280456
rect 118713 280316 118719 280444
rect 118753 280316 118801 280444
rect 118713 280304 118801 280316
rect 117307 280302 117503 280304
rect 117307 280220 117355 280302
rect 117267 280208 117355 280220
rect 115415 280169 115485 280199
rect 114657 280163 114857 280169
rect 114657 280129 114669 280163
rect 114845 280129 114857 280163
rect 114657 280123 114857 280129
rect 115348 280163 115548 280169
rect 115348 280129 115360 280163
rect 115536 280129 115548 280163
rect 115348 280123 115548 280129
rect 112656 279956 112662 280084
rect 112696 279956 112744 280084
rect 113843 280054 114343 280084
rect 113000 280048 114343 280054
rect 113000 280014 113012 280048
rect 114088 280043 114343 280048
rect 114570 280101 114616 280113
rect 114088 280014 114100 280043
rect 113000 280008 114100 280014
rect 112656 279944 112744 279956
rect 111404 279736 111446 279944
rect 111524 279928 112624 279934
rect 111524 279894 111536 279928
rect 112612 279894 112624 279928
rect 111524 279888 112624 279894
rect 111524 279786 112624 279792
rect 111524 279752 111536 279786
rect 112612 279752 112624 279786
rect 111524 279746 112624 279752
rect 112702 279736 112744 279944
rect 111404 279724 111492 279736
rect 111404 279596 111452 279724
rect 111486 279596 111492 279724
rect 111404 279584 111492 279596
rect 112656 279724 112744 279736
rect 112656 279596 112662 279724
rect 112696 279596 112744 279724
rect 112656 279584 112744 279596
rect 112874 279986 112968 279998
rect 112874 279938 112928 279986
rect 112962 279938 112968 279986
rect 112874 279926 112968 279938
rect 114132 279986 114226 279998
rect 114132 279938 114138 279986
rect 114172 279938 114226 279986
rect 114132 279926 114226 279938
rect 112874 279834 112922 279926
rect 113000 279910 114100 279916
rect 113000 279876 113012 279910
rect 114088 279876 114100 279910
rect 113000 279870 114100 279876
rect 114178 279834 114226 279926
rect 112874 279790 114226 279834
rect 114324 279976 114396 279992
rect 114324 279893 114342 279976
rect 114377 279893 114396 279976
rect 114570 279973 114576 280101
rect 114610 279973 114616 280101
rect 114570 279961 114616 279973
rect 114898 280101 114944 280113
rect 114898 279973 114904 280101
rect 114938 279973 114944 280101
rect 114898 279961 114944 279973
rect 115261 280101 115307 280113
rect 115261 279973 115267 280101
rect 115301 279973 115307 280101
rect 115261 279961 115307 279973
rect 115589 280101 115635 280113
rect 115589 279973 115595 280101
rect 115629 279973 115635 280101
rect 115862 280084 115897 280199
rect 116135 280192 117235 280198
rect 116135 280158 116147 280192
rect 117223 280158 117235 280192
rect 116135 280152 117235 280158
rect 117461 280096 117503 280302
rect 117581 280288 118681 280294
rect 117581 280254 117593 280288
rect 118669 280254 118681 280288
rect 117581 280248 118681 280254
rect 117581 280146 118681 280152
rect 117581 280112 117593 280146
rect 118669 280112 118681 280146
rect 117581 280106 118681 280112
rect 118759 280096 118801 280304
rect 117461 280084 117549 280096
rect 115862 280054 116362 280084
rect 115862 280048 117205 280054
rect 115862 280043 116117 280048
rect 116105 280014 116117 280043
rect 117193 280014 117205 280048
rect 116105 280008 117205 280014
rect 115589 279961 115635 279973
rect 115809 279976 115881 279992
rect 114657 279945 114857 279951
rect 114657 279911 114669 279945
rect 114845 279911 114857 279945
rect 114657 279905 114857 279911
rect 115348 279945 115548 279951
rect 115348 279911 115360 279945
rect 115536 279911 115548 279945
rect 115348 279905 115548 279911
rect 114324 279861 114396 279893
rect 115809 279893 115828 279976
rect 115863 279893 115881 279976
rect 114843 279861 115030 279876
rect 114324 279816 114781 279861
rect 112874 279700 112922 279790
rect 113000 279750 114100 279756
rect 113000 279716 113012 279750
rect 114088 279716 114100 279750
rect 113000 279710 114100 279716
rect 114178 279700 114226 279790
rect 114737 279761 114781 279816
rect 114843 279809 114868 279861
rect 114966 279809 115030 279861
rect 114843 279791 115030 279809
rect 115175 279861 115362 279876
rect 115809 279861 115881 279893
rect 115175 279809 115239 279861
rect 115337 279809 115362 279861
rect 115175 279791 115362 279809
rect 115424 279816 115881 279861
rect 115979 279986 116073 279998
rect 115979 279938 116033 279986
rect 116067 279938 116073 279986
rect 115979 279926 116073 279938
rect 117237 279986 117331 279998
rect 117237 279938 117243 279986
rect 117277 279938 117331 279986
rect 117237 279926 117331 279938
rect 115979 279834 116027 279926
rect 116105 279910 117205 279916
rect 116105 279876 116117 279910
rect 117193 279876 117205 279910
rect 116105 279870 117205 279876
rect 117283 279834 117331 279926
rect 115424 279761 115468 279816
rect 115979 279790 117331 279834
rect 114657 279755 114857 279761
rect 114657 279721 114669 279755
rect 114845 279721 114857 279755
rect 114657 279715 114857 279721
rect 115348 279755 115548 279761
rect 115348 279721 115360 279755
rect 115536 279721 115548 279755
rect 115348 279715 115548 279721
rect 112874 279688 112968 279700
rect 112874 279640 112928 279688
rect 112962 279640 112968 279688
rect 112874 279628 112968 279640
rect 114132 279688 114226 279700
rect 114132 279640 114138 279688
rect 114172 279640 114226 279688
rect 114132 279628 114226 279640
rect 114570 279693 114616 279705
rect 111524 279568 112624 279574
rect 111524 279534 111536 279568
rect 112612 279534 112624 279568
rect 111524 279530 112624 279534
rect 112874 279534 112922 279628
rect 114327 279623 114395 279624
rect 114570 279623 114576 279693
rect 113000 279612 114100 279618
rect 113000 279578 113012 279612
rect 114088 279578 114100 279612
rect 113000 279572 114100 279578
rect 114327 279565 114576 279623
rect 114610 279565 114616 279693
rect 114327 279563 114616 279565
rect 114327 279534 114395 279563
rect 114570 279553 114616 279563
rect 114898 279693 114944 279705
rect 114898 279565 114904 279693
rect 114938 279565 114944 279693
rect 114898 279553 114944 279565
rect 115261 279693 115307 279705
rect 115261 279565 115267 279693
rect 115301 279565 115307 279693
rect 115261 279553 115307 279565
rect 115589 279693 115635 279705
rect 115589 279565 115595 279693
rect 115629 279623 115635 279693
rect 115979 279700 116027 279790
rect 116105 279750 117205 279756
rect 116105 279716 116117 279750
rect 117193 279716 117205 279750
rect 116105 279710 117205 279716
rect 117283 279700 117331 279790
rect 115979 279688 116073 279700
rect 115979 279640 116033 279688
rect 116067 279640 116073 279688
rect 115979 279628 116073 279640
rect 117237 279688 117331 279700
rect 117237 279640 117243 279688
rect 117277 279640 117331 279688
rect 117237 279628 117331 279640
rect 115810 279623 115878 279624
rect 115629 279565 115878 279623
rect 116105 279612 117205 279618
rect 116105 279578 116117 279612
rect 117193 279578 117205 279612
rect 116105 279572 117205 279578
rect 115589 279563 115878 279565
rect 115589 279553 115635 279563
rect 112874 279530 114395 279534
rect 111524 279528 114395 279530
rect 112044 279494 114395 279528
rect 114657 279537 114857 279543
rect 114657 279503 114669 279537
rect 114845 279503 114857 279537
rect 114657 279497 114857 279503
rect 115348 279537 115548 279543
rect 115348 279503 115360 279537
rect 115536 279503 115548 279537
rect 115348 279497 115548 279503
rect 115810 279534 115878 279563
rect 117283 279534 117331 279628
rect 117461 279956 117509 280084
rect 117543 279956 117549 280084
rect 117461 279944 117549 279956
rect 118713 280084 118801 280096
rect 118713 279956 118719 280084
rect 118753 279956 118801 280084
rect 118713 279944 118801 279956
rect 117461 279736 117503 279944
rect 117581 279928 118681 279934
rect 117581 279894 117593 279928
rect 118669 279894 118681 279928
rect 117581 279888 118681 279894
rect 117581 279786 118681 279792
rect 117581 279752 117593 279786
rect 118669 279752 118681 279786
rect 117581 279746 118681 279752
rect 118759 279736 118801 279944
rect 117461 279724 117549 279736
rect 117461 279596 117509 279724
rect 117543 279596 117549 279724
rect 117461 279584 117549 279596
rect 118713 279724 118801 279736
rect 118713 279596 118719 279724
rect 118753 279596 118801 279724
rect 118713 279584 118801 279596
rect 115810 279530 117331 279534
rect 117581 279568 118681 279574
rect 117581 279534 117593 279568
rect 118669 279534 118681 279568
rect 117581 279530 118681 279534
rect 115810 279528 118681 279530
rect 112719 279452 112924 279494
rect 113982 279420 114266 279430
rect 114724 279420 114783 279497
rect 113982 279417 114783 279420
rect 113982 279348 114010 279417
rect 114237 279348 114783 279417
rect 113982 279331 114783 279348
rect 115422 279420 115481 279497
rect 115810 279494 118161 279528
rect 117281 279452 117486 279494
rect 115939 279420 116223 279430
rect 115422 279417 116223 279420
rect 115422 279348 115968 279417
rect 116195 279348 116223 279417
rect 115422 279331 116223 279348
rect 113982 279330 114266 279331
rect 115939 279330 116223 279331
rect 112970 279208 114070 279214
rect 111524 279200 112624 279206
rect 111524 279166 111536 279200
rect 112612 279166 112624 279200
rect 112970 279174 112982 279208
rect 114058 279174 114070 279208
rect 116135 279208 117235 279214
rect 112970 279168 114070 279174
rect 114657 279183 114857 279189
rect 111524 279160 112624 279166
rect 111404 279138 111492 279150
rect 111404 279010 111452 279138
rect 111486 279010 111492 279138
rect 111404 278998 111492 279010
rect 112656 279138 112744 279150
rect 112656 279010 112662 279138
rect 112696 279082 112744 279138
rect 112850 279146 112938 279158
rect 112850 279082 112898 279146
rect 112696 279020 112898 279082
rect 112696 279010 112744 279020
rect 112656 278998 112744 279010
rect 111404 278790 111446 278998
rect 111524 278982 112624 278988
rect 111524 278948 111536 278982
rect 112612 278948 112624 278982
rect 111524 278942 112624 278948
rect 112702 278966 112744 278998
rect 112850 278978 112898 279020
rect 112932 278978 112938 279146
rect 112850 278966 112938 278978
rect 114102 279146 114190 279158
rect 114102 278978 114108 279146
rect 114142 279092 114190 279146
rect 114657 279149 114669 279183
rect 114845 279149 114857 279183
rect 114657 279143 114857 279149
rect 115348 279183 115548 279189
rect 115348 279149 115360 279183
rect 115536 279149 115548 279183
rect 116135 279174 116147 279208
rect 117223 279174 117235 279208
rect 116135 279168 117235 279174
rect 117581 279200 118681 279206
rect 117581 279166 117593 279200
rect 118669 279166 118681 279200
rect 117581 279160 118681 279166
rect 115348 279143 115548 279149
rect 116015 279146 116103 279158
rect 114570 279121 114616 279133
rect 114570 279092 114576 279121
rect 114142 278978 114576 279092
rect 114102 278966 114576 278978
rect 111524 278840 112624 278846
rect 111524 278806 111536 278840
rect 112612 278806 112624 278840
rect 111524 278800 112624 278806
rect 112702 278790 112746 278966
rect 111404 278778 111492 278790
rect 111404 278650 111452 278778
rect 111486 278650 111492 278778
rect 111404 278638 111492 278650
rect 112656 278778 112746 278790
rect 112656 278650 112662 278778
rect 112696 278746 112746 278778
rect 112850 278866 112892 278966
rect 114148 278959 114576 278966
rect 112970 278950 114070 278956
rect 112970 278916 112982 278950
rect 114058 278916 114070 278950
rect 112970 278910 114070 278916
rect 114148 278866 114190 278959
rect 112850 278828 114190 278866
rect 112696 278698 112744 278746
rect 112850 278734 112892 278828
rect 112970 278784 114070 278790
rect 112970 278750 112982 278784
rect 114058 278750 114070 278784
rect 112970 278744 114070 278750
rect 114148 278734 114190 278828
rect 114570 278753 114576 278959
rect 114610 278753 114616 279121
rect 114570 278741 114616 278753
rect 114898 279121 114944 279133
rect 114898 278753 114904 279121
rect 114938 278753 114944 279121
rect 114898 278741 114944 278753
rect 115261 279121 115307 279133
rect 115261 278753 115267 279121
rect 115301 278753 115307 279121
rect 115261 278741 115307 278753
rect 115589 279121 115635 279133
rect 115589 278753 115595 279121
rect 115629 279092 115635 279121
rect 116015 279092 116063 279146
rect 115629 278978 116063 279092
rect 116097 278978 116103 279146
rect 115629 278966 116103 278978
rect 117267 279146 117355 279158
rect 117267 278978 117273 279146
rect 117307 279082 117355 279146
rect 117461 279138 117549 279150
rect 117461 279082 117509 279138
rect 117307 279020 117509 279082
rect 117307 278978 117355 279020
rect 117267 278966 117355 278978
rect 117461 279010 117509 279020
rect 117543 279010 117549 279138
rect 117461 278998 117549 279010
rect 118713 279138 118801 279150
rect 118713 279010 118719 279138
rect 118753 279010 118801 279138
rect 118713 278998 118801 279010
rect 117461 278966 117503 278998
rect 115629 278959 116057 278966
rect 115629 278753 115635 278959
rect 115589 278741 115635 278753
rect 116015 278866 116057 278959
rect 116135 278950 117235 278956
rect 116135 278916 116147 278950
rect 117223 278916 117235 278950
rect 116135 278910 117235 278916
rect 117313 278866 117355 278966
rect 116015 278828 117355 278866
rect 112850 278722 112938 278734
rect 112850 278698 112898 278722
rect 112696 278650 112898 278698
rect 112656 278638 112898 278650
rect 111404 278430 111446 278638
rect 112702 278636 112898 278638
rect 111524 278622 112624 278628
rect 111524 278588 111536 278622
rect 112612 278588 112624 278622
rect 111524 278582 112624 278588
rect 111524 278480 112624 278486
rect 111524 278446 111536 278480
rect 112612 278446 112624 278480
rect 111524 278440 112624 278446
rect 112702 278430 112744 278636
rect 112850 278554 112898 278636
rect 112932 278554 112938 278722
rect 112850 278542 112938 278554
rect 114102 278722 114190 278734
rect 116015 278734 116057 278828
rect 116135 278784 117235 278790
rect 116135 278750 116147 278784
rect 117223 278750 117235 278784
rect 116135 278744 117235 278750
rect 117313 278734 117355 278828
rect 117459 278790 117503 278966
rect 117581 278982 118681 278988
rect 117581 278948 117593 278982
rect 118669 278948 118681 278982
rect 117581 278942 118681 278948
rect 117581 278840 118681 278846
rect 117581 278806 117593 278840
rect 118669 278806 118681 278840
rect 117581 278800 118681 278806
rect 118759 278790 118801 278998
rect 117459 278778 117549 278790
rect 117459 278746 117509 278778
rect 114102 278554 114108 278722
rect 114142 278554 114190 278722
rect 114657 278725 114857 278731
rect 114657 278691 114669 278725
rect 114845 278691 114857 278725
rect 114657 278685 114857 278691
rect 115348 278725 115548 278731
rect 115348 278691 115360 278725
rect 115536 278691 115548 278725
rect 115348 278685 115548 278691
rect 116015 278722 116103 278734
rect 114720 278617 114790 278685
rect 114102 278542 114190 278554
rect 114308 278533 114790 278617
rect 114865 278628 114970 278645
rect 114865 278560 114885 278628
rect 114948 278560 114970 278628
rect 114865 278538 114970 278560
rect 115235 278628 115340 278645
rect 115235 278560 115257 278628
rect 115320 278560 115340 278628
rect 115235 278538 115340 278560
rect 115415 278617 115485 278685
rect 112970 278526 114070 278532
rect 112970 278492 112982 278526
rect 114058 278492 114070 278526
rect 112970 278486 114070 278492
rect 111404 278418 111492 278430
rect 111404 278290 111452 278418
rect 111486 278290 111492 278418
rect 111404 278278 111492 278290
rect 112656 278418 112744 278430
rect 114308 278418 114343 278533
rect 114720 278503 114790 278533
rect 115415 278533 115897 278617
rect 116015 278554 116063 278722
rect 116097 278554 116103 278722
rect 116015 278542 116103 278554
rect 117267 278722 117355 278734
rect 117267 278554 117273 278722
rect 117307 278698 117355 278722
rect 117461 278698 117509 278746
rect 117307 278650 117509 278698
rect 117543 278650 117549 278778
rect 117307 278638 117549 278650
rect 118713 278778 118801 278790
rect 118713 278650 118719 278778
rect 118753 278650 118801 278778
rect 118713 278638 118801 278650
rect 117307 278636 117503 278638
rect 117307 278554 117355 278636
rect 117267 278542 117355 278554
rect 115415 278503 115485 278533
rect 114657 278497 114857 278503
rect 114657 278463 114669 278497
rect 114845 278463 114857 278497
rect 114657 278457 114857 278463
rect 115348 278497 115548 278503
rect 115348 278463 115360 278497
rect 115536 278463 115548 278497
rect 115348 278457 115548 278463
rect 112656 278290 112662 278418
rect 112696 278290 112744 278418
rect 113843 278388 114343 278418
rect 113000 278382 114343 278388
rect 113000 278348 113012 278382
rect 114088 278377 114343 278382
rect 114570 278435 114616 278447
rect 114088 278348 114100 278377
rect 113000 278342 114100 278348
rect 112656 278278 112744 278290
rect 111404 278070 111446 278278
rect 111524 278262 112624 278268
rect 111524 278228 111536 278262
rect 112612 278228 112624 278262
rect 111524 278222 112624 278228
rect 111524 278120 112624 278126
rect 111524 278086 111536 278120
rect 112612 278086 112624 278120
rect 111524 278080 112624 278086
rect 112702 278070 112744 278278
rect 111404 278058 111492 278070
rect 111404 277930 111452 278058
rect 111486 277930 111492 278058
rect 111404 277918 111492 277930
rect 112656 278058 112744 278070
rect 112656 277930 112662 278058
rect 112696 277930 112744 278058
rect 112656 277918 112744 277930
rect 112874 278320 112968 278332
rect 112874 278272 112928 278320
rect 112962 278272 112968 278320
rect 112874 278260 112968 278272
rect 114132 278320 114226 278332
rect 114132 278272 114138 278320
rect 114172 278272 114226 278320
rect 114132 278260 114226 278272
rect 112874 278168 112922 278260
rect 113000 278244 114100 278250
rect 113000 278210 113012 278244
rect 114088 278210 114100 278244
rect 113000 278204 114100 278210
rect 114178 278168 114226 278260
rect 112874 278124 114226 278168
rect 114324 278310 114396 278326
rect 114324 278227 114342 278310
rect 114377 278227 114396 278310
rect 114570 278307 114576 278435
rect 114610 278307 114616 278435
rect 114570 278295 114616 278307
rect 114898 278435 114944 278447
rect 114898 278307 114904 278435
rect 114938 278307 114944 278435
rect 114898 278295 114944 278307
rect 115261 278435 115307 278447
rect 115261 278307 115267 278435
rect 115301 278307 115307 278435
rect 115261 278295 115307 278307
rect 115589 278435 115635 278447
rect 115589 278307 115595 278435
rect 115629 278307 115635 278435
rect 115862 278418 115897 278533
rect 116135 278526 117235 278532
rect 116135 278492 116147 278526
rect 117223 278492 117235 278526
rect 116135 278486 117235 278492
rect 117461 278430 117503 278636
rect 117581 278622 118681 278628
rect 117581 278588 117593 278622
rect 118669 278588 118681 278622
rect 117581 278582 118681 278588
rect 117581 278480 118681 278486
rect 117581 278446 117593 278480
rect 118669 278446 118681 278480
rect 117581 278440 118681 278446
rect 118759 278430 118801 278638
rect 119257 278715 119341 281145
rect 119757 278715 119845 281145
rect 124495 280818 124958 280846
rect 123506 280816 124958 280818
rect 123444 280811 124958 280816
rect 121846 280796 124958 280811
rect 120433 280718 120825 280724
rect 120433 280684 120445 280718
rect 120813 280684 120825 280718
rect 120433 280678 120825 280684
rect 121133 280718 121525 280724
rect 121133 280684 121145 280718
rect 121513 280684 121525 280718
rect 121133 280678 121525 280684
rect 121846 280696 124552 280796
rect 120377 280625 120423 280637
rect 120377 280549 120383 280625
rect 120417 280549 120423 280625
rect 120377 280537 120423 280549
rect 120835 280625 120881 280637
rect 120835 280549 120841 280625
rect 120875 280549 120881 280625
rect 120835 280537 120881 280549
rect 121077 280625 121123 280637
rect 121077 280549 121083 280625
rect 121117 280549 121123 280625
rect 121077 280537 121123 280549
rect 121535 280625 121581 280637
rect 121535 280549 121541 280625
rect 121575 280549 121581 280625
rect 121535 280537 121581 280549
rect 120433 280490 120825 280496
rect 120433 280456 120445 280490
rect 120813 280456 120825 280490
rect 120433 280450 120825 280456
rect 121133 280490 121525 280496
rect 121133 280456 121145 280490
rect 121513 280456 121525 280490
rect 121133 280450 121525 280456
rect 121846 280383 121915 280696
rect 123444 280632 124552 280696
rect 123444 280510 123545 280632
rect 124495 280559 124552 280632
rect 124902 280559 124958 280796
rect 122360 280504 122752 280510
rect 122360 280470 122372 280504
rect 122740 280470 122752 280504
rect 122360 280464 122752 280470
rect 123060 280504 123551 280510
rect 123060 280470 123072 280504
rect 123440 280470 123551 280504
rect 124495 280498 124958 280559
rect 123060 280464 123551 280470
rect 123452 280423 123551 280464
rect 121134 280340 121915 280383
rect 120433 280334 120825 280340
rect 120433 280300 120445 280334
rect 120813 280300 120825 280334
rect 120433 280294 120825 280300
rect 121133 280339 121915 280340
rect 122304 280411 122350 280423
rect 121133 280334 121525 280339
rect 121133 280300 121145 280334
rect 121513 280300 121525 280334
rect 121133 280294 121525 280300
rect 120377 280241 120423 280253
rect 120377 279765 120383 280241
rect 120417 279765 120423 280241
rect 120377 279753 120423 279765
rect 120835 280241 120881 280253
rect 120835 279765 120841 280241
rect 120875 280064 120881 280241
rect 121077 280241 121123 280253
rect 121077 280064 121083 280241
rect 120875 279937 121083 280064
rect 120875 279765 120881 279937
rect 120835 279753 120881 279765
rect 120433 279706 120825 279712
rect 120433 279672 120445 279706
rect 120813 279672 120825 279706
rect 120433 279656 120825 279672
rect 120433 279564 120501 279656
rect 120737 279564 120825 279656
rect 120433 279550 120825 279564
rect 120433 279516 120445 279550
rect 120813 279516 120825 279550
rect 120433 279510 120825 279516
rect 120377 279457 120423 279469
rect 120377 278981 120383 279457
rect 120417 278981 120423 279457
rect 120377 278969 120423 278981
rect 120835 279457 120881 279469
rect 120835 278981 120841 279457
rect 120875 279280 120881 279457
rect 120953 279280 121018 279937
rect 121077 279765 121083 279937
rect 121117 279765 121123 280241
rect 121077 279753 121123 279765
rect 121535 280241 121624 280253
rect 121535 279765 121541 280241
rect 121575 279765 121624 280241
rect 121535 279753 121624 279765
rect 121133 279706 121525 279712
rect 121133 279672 121145 279706
rect 121513 279672 121525 279706
rect 121133 279550 121525 279672
rect 121133 279516 121145 279550
rect 121513 279516 121525 279550
rect 121133 279510 121525 279516
rect 121581 279469 121624 279753
rect 121797 279887 122235 279937
rect 122304 279935 122310 280411
rect 122344 279935 122350 280411
rect 122304 279923 122350 279935
rect 122762 280411 123050 280423
rect 122762 279935 122768 280411
rect 122802 279935 123010 280411
rect 123044 279935 123050 280411
rect 122762 279923 123050 279935
rect 123462 280411 123551 280423
rect 123462 279935 123468 280411
rect 123502 279935 123551 280411
rect 123462 279923 123551 279935
rect 121077 279457 121123 279469
rect 121077 279280 121083 279457
rect 120875 279153 121083 279280
rect 120875 278981 120881 279153
rect 120835 278969 120881 278981
rect 120433 278922 120825 278928
rect 120433 278888 120445 278922
rect 120813 278888 120825 278922
rect 120433 278766 120825 278888
rect 120433 278732 120445 278766
rect 120813 278732 120825 278766
rect 120433 278726 120825 278732
rect 119257 278619 119845 278715
rect 120377 278673 120423 278685
rect 117461 278418 117549 278430
rect 115862 278388 116362 278418
rect 115862 278382 117205 278388
rect 115862 278377 116117 278382
rect 116105 278348 116117 278377
rect 117193 278348 117205 278382
rect 116105 278342 117205 278348
rect 115589 278295 115635 278307
rect 115809 278310 115881 278326
rect 114657 278279 114857 278285
rect 114657 278245 114669 278279
rect 114845 278245 114857 278279
rect 114657 278239 114857 278245
rect 115348 278279 115548 278285
rect 115348 278245 115360 278279
rect 115536 278245 115548 278279
rect 115348 278239 115548 278245
rect 114324 278195 114396 278227
rect 115809 278227 115828 278310
rect 115863 278227 115881 278310
rect 114843 278195 115030 278210
rect 114324 278150 114781 278195
rect 112874 278034 112922 278124
rect 113000 278084 114100 278090
rect 113000 278050 113012 278084
rect 114088 278050 114100 278084
rect 113000 278044 114100 278050
rect 114178 278034 114226 278124
rect 114737 278095 114781 278150
rect 114843 278143 114868 278195
rect 114966 278143 115030 278195
rect 114843 278125 115030 278143
rect 115175 278195 115362 278210
rect 115809 278195 115881 278227
rect 115175 278143 115239 278195
rect 115337 278143 115362 278195
rect 115175 278125 115362 278143
rect 115424 278150 115881 278195
rect 115979 278320 116073 278332
rect 115979 278272 116033 278320
rect 116067 278272 116073 278320
rect 115979 278260 116073 278272
rect 117237 278320 117331 278332
rect 117237 278272 117243 278320
rect 117277 278272 117331 278320
rect 117237 278260 117331 278272
rect 115979 278168 116027 278260
rect 116105 278244 117205 278250
rect 116105 278210 116117 278244
rect 117193 278210 117205 278244
rect 116105 278204 117205 278210
rect 117283 278168 117331 278260
rect 115424 278095 115468 278150
rect 115979 278124 117331 278168
rect 114657 278089 114857 278095
rect 114657 278055 114669 278089
rect 114845 278055 114857 278089
rect 114657 278049 114857 278055
rect 115348 278089 115548 278095
rect 115348 278055 115360 278089
rect 115536 278055 115548 278089
rect 115348 278049 115548 278055
rect 112874 278022 112968 278034
rect 112874 277974 112928 278022
rect 112962 277974 112968 278022
rect 112874 277962 112968 277974
rect 114132 278022 114226 278034
rect 114132 277974 114138 278022
rect 114172 277974 114226 278022
rect 114132 277962 114226 277974
rect 114570 278027 114616 278039
rect 111524 277902 112624 277908
rect 111524 277868 111536 277902
rect 112612 277868 112624 277902
rect 111524 277864 112624 277868
rect 112874 277868 112922 277962
rect 114327 277957 114395 277958
rect 114570 277957 114576 278027
rect 113000 277946 114100 277952
rect 113000 277912 113012 277946
rect 114088 277912 114100 277946
rect 113000 277906 114100 277912
rect 114327 277899 114576 277957
rect 114610 277899 114616 278027
rect 114327 277897 114616 277899
rect 114327 277868 114395 277897
rect 114570 277887 114616 277897
rect 114898 278027 114944 278039
rect 114898 277899 114904 278027
rect 114938 277899 114944 278027
rect 114898 277887 114944 277899
rect 115261 278027 115307 278039
rect 115261 277899 115267 278027
rect 115301 277899 115307 278027
rect 115261 277887 115307 277899
rect 115589 278027 115635 278039
rect 115589 277899 115595 278027
rect 115629 277957 115635 278027
rect 115979 278034 116027 278124
rect 116105 278084 117205 278090
rect 116105 278050 116117 278084
rect 117193 278050 117205 278084
rect 116105 278044 117205 278050
rect 117283 278034 117331 278124
rect 115979 278022 116073 278034
rect 115979 277974 116033 278022
rect 116067 277974 116073 278022
rect 115979 277962 116073 277974
rect 117237 278022 117331 278034
rect 117237 277974 117243 278022
rect 117277 277974 117331 278022
rect 117237 277962 117331 277974
rect 115810 277957 115878 277958
rect 115629 277899 115878 277957
rect 116105 277946 117205 277952
rect 116105 277912 116117 277946
rect 117193 277912 117205 277946
rect 116105 277906 117205 277912
rect 115589 277897 115878 277899
rect 115589 277887 115635 277897
rect 112874 277864 114395 277868
rect 111524 277862 114395 277864
rect 112044 277828 114395 277862
rect 114657 277871 114857 277877
rect 114657 277837 114669 277871
rect 114845 277837 114857 277871
rect 114657 277831 114857 277837
rect 115348 277871 115548 277877
rect 115348 277837 115360 277871
rect 115536 277837 115548 277871
rect 115348 277831 115548 277837
rect 115810 277868 115878 277897
rect 117283 277868 117331 277962
rect 117461 278290 117509 278418
rect 117543 278290 117549 278418
rect 117461 278278 117549 278290
rect 118713 278418 118801 278430
rect 118713 278290 118719 278418
rect 118753 278290 118801 278418
rect 118713 278278 118801 278290
rect 117461 278070 117503 278278
rect 117581 278262 118681 278268
rect 117581 278228 117593 278262
rect 118669 278228 118681 278262
rect 117581 278222 118681 278228
rect 117581 278120 118681 278126
rect 117581 278086 117593 278120
rect 118669 278086 118681 278120
rect 117581 278080 118681 278086
rect 118759 278070 118801 278278
rect 120377 278197 120383 278673
rect 120417 278197 120423 278673
rect 120377 278185 120423 278197
rect 120835 278673 120881 278685
rect 120835 278197 120841 278673
rect 120875 278496 120881 278673
rect 120953 278496 121018 279153
rect 121077 278981 121083 279153
rect 121117 278981 121123 279457
rect 121077 278969 121123 278981
rect 121535 279457 121677 279469
rect 121535 278981 121541 279457
rect 121575 279396 121677 279457
rect 121575 278981 121605 279396
rect 121535 278969 121605 278981
rect 121133 278922 121525 278928
rect 121133 278888 121145 278922
rect 121513 278888 121525 278922
rect 121133 278766 121525 278888
rect 121133 278732 121145 278766
rect 121513 278732 121525 278766
rect 121133 278726 121525 278732
rect 121581 278685 121605 278969
rect 121077 278673 121123 278685
rect 121077 278496 121083 278673
rect 120875 278369 121083 278496
rect 120875 278197 120881 278369
rect 120835 278185 120881 278197
rect 117461 278058 117549 278070
rect 117461 277930 117509 278058
rect 117543 277930 117549 278058
rect 117461 277918 117549 277930
rect 118713 278058 118801 278070
rect 118713 277930 118719 278058
rect 118753 277930 118801 278058
rect 120433 278138 120825 278144
rect 120433 278104 120445 278138
rect 120813 278104 120825 278138
rect 120433 277982 120825 278104
rect 120433 277948 120445 277982
rect 120813 277948 120825 277982
rect 120433 277942 120825 277948
rect 118713 277918 118801 277930
rect 115810 277864 117331 277868
rect 117581 277902 118681 277908
rect 117581 277868 117593 277902
rect 118669 277868 118681 277902
rect 117581 277864 118681 277868
rect 115810 277862 118681 277864
rect 120377 277889 120423 277901
rect 112719 277786 112924 277828
rect 113982 277754 114266 277764
rect 114724 277754 114783 277831
rect 113982 277751 114783 277754
rect 113982 277682 114010 277751
rect 114237 277682 114783 277751
rect 113982 277665 114783 277682
rect 115422 277754 115481 277831
rect 115810 277828 118161 277862
rect 117281 277786 117486 277828
rect 115939 277754 116223 277764
rect 115422 277751 116223 277754
rect 115422 277682 115968 277751
rect 116195 277682 116223 277751
rect 115422 277665 116223 277682
rect 113982 277664 114266 277665
rect 115939 277664 116223 277665
rect 112970 277542 114070 277548
rect 111524 277534 112624 277540
rect 111524 277500 111536 277534
rect 112612 277500 112624 277534
rect 112970 277508 112982 277542
rect 114058 277508 114070 277542
rect 116135 277542 117235 277548
rect 112970 277502 114070 277508
rect 114657 277517 114857 277523
rect 111524 277494 112624 277500
rect 111404 277472 111492 277484
rect 111404 277344 111452 277472
rect 111486 277344 111492 277472
rect 111404 277332 111492 277344
rect 112656 277472 112744 277484
rect 112656 277344 112662 277472
rect 112696 277416 112744 277472
rect 112850 277480 112938 277492
rect 112850 277416 112898 277480
rect 112696 277354 112898 277416
rect 112696 277344 112744 277354
rect 112656 277332 112744 277344
rect 111404 277124 111446 277332
rect 111524 277316 112624 277322
rect 111524 277282 111536 277316
rect 112612 277282 112624 277316
rect 111524 277276 112624 277282
rect 112702 277300 112744 277332
rect 112850 277312 112898 277354
rect 112932 277312 112938 277480
rect 112850 277300 112938 277312
rect 114102 277480 114190 277492
rect 114102 277312 114108 277480
rect 114142 277426 114190 277480
rect 114657 277483 114669 277517
rect 114845 277483 114857 277517
rect 114657 277477 114857 277483
rect 115348 277517 115548 277523
rect 115348 277483 115360 277517
rect 115536 277483 115548 277517
rect 116135 277508 116147 277542
rect 117223 277508 117235 277542
rect 116135 277502 117235 277508
rect 117581 277534 118681 277540
rect 117581 277500 117593 277534
rect 118669 277500 118681 277534
rect 117581 277494 118681 277500
rect 115348 277477 115548 277483
rect 116015 277480 116103 277492
rect 114570 277455 114616 277467
rect 114570 277426 114576 277455
rect 114142 277312 114576 277426
rect 114102 277300 114576 277312
rect 111524 277174 112624 277180
rect 111524 277140 111536 277174
rect 112612 277140 112624 277174
rect 111524 277134 112624 277140
rect 112702 277124 112746 277300
rect 111404 277112 111492 277124
rect 111404 276984 111452 277112
rect 111486 276984 111492 277112
rect 111404 276972 111492 276984
rect 112656 277112 112746 277124
rect 112656 276984 112662 277112
rect 112696 277080 112746 277112
rect 112850 277200 112892 277300
rect 114148 277293 114576 277300
rect 112970 277284 114070 277290
rect 112970 277250 112982 277284
rect 114058 277250 114070 277284
rect 112970 277244 114070 277250
rect 114148 277200 114190 277293
rect 112850 277162 114190 277200
rect 112696 277032 112744 277080
rect 112850 277068 112892 277162
rect 112970 277118 114070 277124
rect 112970 277084 112982 277118
rect 114058 277084 114070 277118
rect 112970 277078 114070 277084
rect 114148 277068 114190 277162
rect 114570 277087 114576 277293
rect 114610 277087 114616 277455
rect 114570 277075 114616 277087
rect 114898 277455 114944 277467
rect 114898 277087 114904 277455
rect 114938 277087 114944 277455
rect 114898 277075 114944 277087
rect 115261 277455 115307 277467
rect 115261 277087 115267 277455
rect 115301 277087 115307 277455
rect 115261 277075 115307 277087
rect 115589 277455 115635 277467
rect 115589 277087 115595 277455
rect 115629 277426 115635 277455
rect 116015 277426 116063 277480
rect 115629 277312 116063 277426
rect 116097 277312 116103 277480
rect 115629 277300 116103 277312
rect 117267 277480 117355 277492
rect 117267 277312 117273 277480
rect 117307 277416 117355 277480
rect 117461 277472 117549 277484
rect 117461 277416 117509 277472
rect 117307 277354 117509 277416
rect 117307 277312 117355 277354
rect 117267 277300 117355 277312
rect 117461 277344 117509 277354
rect 117543 277344 117549 277472
rect 117461 277332 117549 277344
rect 118713 277472 118801 277484
rect 118713 277344 118719 277472
rect 118753 277344 118801 277472
rect 120377 277413 120383 277889
rect 120417 277413 120423 277889
rect 120377 277401 120423 277413
rect 120835 277889 120881 277901
rect 120835 277413 120841 277889
rect 120875 277712 120881 277889
rect 120953 277712 121018 278369
rect 121077 278197 121083 278369
rect 121117 278197 121123 278673
rect 121077 278185 121123 278197
rect 121535 278673 121605 278685
rect 121535 278197 121541 278673
rect 121575 278197 121605 278673
rect 121535 278185 121605 278197
rect 121133 278138 121525 278144
rect 121133 278104 121145 278138
rect 121513 278104 121525 278138
rect 121133 277982 121525 278104
rect 121133 277948 121145 277982
rect 121513 277948 121525 277982
rect 121133 277942 121525 277948
rect 121581 277901 121605 278185
rect 121077 277889 121123 277901
rect 121077 277712 121083 277889
rect 120875 277585 121083 277712
rect 120875 277413 120881 277585
rect 120835 277401 120881 277413
rect 118713 277332 118801 277344
rect 117461 277300 117503 277332
rect 115629 277293 116057 277300
rect 115629 277087 115635 277293
rect 115589 277075 115635 277087
rect 116015 277200 116057 277293
rect 116135 277284 117235 277290
rect 116135 277250 116147 277284
rect 117223 277250 117235 277284
rect 116135 277244 117235 277250
rect 117313 277200 117355 277300
rect 116015 277162 117355 277200
rect 112850 277056 112938 277068
rect 112850 277032 112898 277056
rect 112696 276984 112898 277032
rect 112656 276972 112898 276984
rect 111404 276764 111446 276972
rect 112702 276970 112898 276972
rect 111524 276956 112624 276962
rect 111524 276922 111536 276956
rect 112612 276922 112624 276956
rect 111524 276916 112624 276922
rect 111524 276814 112624 276820
rect 111524 276780 111536 276814
rect 112612 276780 112624 276814
rect 111524 276774 112624 276780
rect 112702 276764 112744 276970
rect 112850 276888 112898 276970
rect 112932 276888 112938 277056
rect 112850 276876 112938 276888
rect 114102 277056 114190 277068
rect 116015 277068 116057 277162
rect 116135 277118 117235 277124
rect 116135 277084 116147 277118
rect 117223 277084 117235 277118
rect 116135 277078 117235 277084
rect 117313 277068 117355 277162
rect 117459 277124 117503 277300
rect 117581 277316 118681 277322
rect 117581 277282 117593 277316
rect 118669 277282 118681 277316
rect 117581 277276 118681 277282
rect 117581 277174 118681 277180
rect 117581 277140 117593 277174
rect 118669 277140 118681 277174
rect 117581 277134 118681 277140
rect 118759 277124 118801 277332
rect 120433 277354 120825 277360
rect 120433 277320 120445 277354
rect 120813 277320 120825 277354
rect 120433 277198 120825 277320
rect 120433 277164 120445 277198
rect 120813 277164 120825 277198
rect 120433 277158 120825 277164
rect 117459 277112 117549 277124
rect 117459 277080 117509 277112
rect 114102 276888 114108 277056
rect 114142 276888 114190 277056
rect 114657 277059 114857 277065
rect 114657 277025 114669 277059
rect 114845 277025 114857 277059
rect 114657 277019 114857 277025
rect 115348 277059 115548 277065
rect 115348 277025 115360 277059
rect 115536 277025 115548 277059
rect 115348 277019 115548 277025
rect 116015 277056 116103 277068
rect 114720 276951 114790 277019
rect 114102 276876 114190 276888
rect 114308 276867 114790 276951
rect 114865 276962 114970 276979
rect 114865 276894 114885 276962
rect 114948 276894 114970 276962
rect 114865 276872 114970 276894
rect 115235 276962 115340 276979
rect 115235 276894 115257 276962
rect 115320 276894 115340 276962
rect 115235 276872 115340 276894
rect 115415 276951 115485 277019
rect 112970 276860 114070 276866
rect 112970 276826 112982 276860
rect 114058 276826 114070 276860
rect 112970 276820 114070 276826
rect 111404 276752 111492 276764
rect 111404 276624 111452 276752
rect 111486 276624 111492 276752
rect 111404 276612 111492 276624
rect 112656 276752 112744 276764
rect 114308 276752 114343 276867
rect 114720 276837 114790 276867
rect 115415 276867 115897 276951
rect 116015 276888 116063 277056
rect 116097 276888 116103 277056
rect 116015 276876 116103 276888
rect 117267 277056 117355 277068
rect 117267 276888 117273 277056
rect 117307 277032 117355 277056
rect 117461 277032 117509 277080
rect 117307 276984 117509 277032
rect 117543 276984 117549 277112
rect 117307 276972 117549 276984
rect 118713 277112 118801 277124
rect 118713 276984 118719 277112
rect 118753 276984 118801 277112
rect 118713 276972 118801 276984
rect 117307 276970 117503 276972
rect 117307 276888 117355 276970
rect 117267 276876 117355 276888
rect 115415 276837 115485 276867
rect 114657 276831 114857 276837
rect 114657 276797 114669 276831
rect 114845 276797 114857 276831
rect 114657 276791 114857 276797
rect 115348 276831 115548 276837
rect 115348 276797 115360 276831
rect 115536 276797 115548 276831
rect 115348 276791 115548 276797
rect 112656 276624 112662 276752
rect 112696 276624 112744 276752
rect 113843 276722 114343 276752
rect 113000 276716 114343 276722
rect 113000 276682 113012 276716
rect 114088 276711 114343 276716
rect 114570 276769 114616 276781
rect 114088 276682 114100 276711
rect 113000 276676 114100 276682
rect 112656 276612 112744 276624
rect 111404 276404 111446 276612
rect 111524 276596 112624 276602
rect 111524 276562 111536 276596
rect 112612 276562 112624 276596
rect 111524 276556 112624 276562
rect 111524 276454 112624 276460
rect 111524 276420 111536 276454
rect 112612 276420 112624 276454
rect 111524 276414 112624 276420
rect 112702 276404 112744 276612
rect 111404 276392 111492 276404
rect 111404 276264 111452 276392
rect 111486 276264 111492 276392
rect 111404 276252 111492 276264
rect 112656 276392 112744 276404
rect 112656 276264 112662 276392
rect 112696 276264 112744 276392
rect 112656 276252 112744 276264
rect 112874 276654 112968 276666
rect 112874 276606 112928 276654
rect 112962 276606 112968 276654
rect 112874 276594 112968 276606
rect 114132 276654 114226 276666
rect 114132 276606 114138 276654
rect 114172 276606 114226 276654
rect 114132 276594 114226 276606
rect 112874 276502 112922 276594
rect 113000 276578 114100 276584
rect 113000 276544 113012 276578
rect 114088 276544 114100 276578
rect 113000 276538 114100 276544
rect 114178 276502 114226 276594
rect 112874 276458 114226 276502
rect 114324 276644 114396 276660
rect 114324 276561 114342 276644
rect 114377 276561 114396 276644
rect 114570 276641 114576 276769
rect 114610 276641 114616 276769
rect 114570 276629 114616 276641
rect 114898 276769 114944 276781
rect 114898 276641 114904 276769
rect 114938 276641 114944 276769
rect 114898 276629 114944 276641
rect 115261 276769 115307 276781
rect 115261 276641 115267 276769
rect 115301 276641 115307 276769
rect 115261 276629 115307 276641
rect 115589 276769 115635 276781
rect 115589 276641 115595 276769
rect 115629 276641 115635 276769
rect 115862 276752 115897 276867
rect 116135 276860 117235 276866
rect 116135 276826 116147 276860
rect 117223 276826 117235 276860
rect 116135 276820 117235 276826
rect 117461 276764 117503 276970
rect 117581 276956 118681 276962
rect 117581 276922 117593 276956
rect 118669 276922 118681 276956
rect 117581 276916 118681 276922
rect 117581 276814 118681 276820
rect 117581 276780 117593 276814
rect 118669 276780 118681 276814
rect 117581 276774 118681 276780
rect 118759 276764 118801 276972
rect 117461 276752 117549 276764
rect 115862 276722 116362 276752
rect 115862 276716 117205 276722
rect 115862 276711 116117 276716
rect 116105 276682 116117 276711
rect 117193 276682 117205 276716
rect 116105 276676 117205 276682
rect 115589 276629 115635 276641
rect 115809 276644 115881 276660
rect 114657 276613 114857 276619
rect 114657 276579 114669 276613
rect 114845 276579 114857 276613
rect 114657 276573 114857 276579
rect 115348 276613 115548 276619
rect 115348 276579 115360 276613
rect 115536 276579 115548 276613
rect 115348 276573 115548 276579
rect 114324 276529 114396 276561
rect 115809 276561 115828 276644
rect 115863 276561 115881 276644
rect 114843 276529 115030 276544
rect 114324 276484 114781 276529
rect 112874 276368 112922 276458
rect 113000 276418 114100 276424
rect 113000 276384 113012 276418
rect 114088 276384 114100 276418
rect 113000 276378 114100 276384
rect 114178 276368 114226 276458
rect 114737 276429 114781 276484
rect 114843 276477 114868 276529
rect 114966 276477 115030 276529
rect 114843 276459 115030 276477
rect 115175 276529 115362 276544
rect 115809 276529 115881 276561
rect 115175 276477 115239 276529
rect 115337 276477 115362 276529
rect 115175 276459 115362 276477
rect 115424 276484 115881 276529
rect 115979 276654 116073 276666
rect 115979 276606 116033 276654
rect 116067 276606 116073 276654
rect 115979 276594 116073 276606
rect 117237 276654 117331 276666
rect 117237 276606 117243 276654
rect 117277 276606 117331 276654
rect 117237 276594 117331 276606
rect 115979 276502 116027 276594
rect 116105 276578 117205 276584
rect 116105 276544 116117 276578
rect 117193 276544 117205 276578
rect 116105 276538 117205 276544
rect 117283 276502 117331 276594
rect 115424 276429 115468 276484
rect 115979 276458 117331 276502
rect 114657 276423 114857 276429
rect 114657 276389 114669 276423
rect 114845 276389 114857 276423
rect 114657 276383 114857 276389
rect 115348 276423 115548 276429
rect 115348 276389 115360 276423
rect 115536 276389 115548 276423
rect 115348 276383 115548 276389
rect 112874 276356 112968 276368
rect 112874 276308 112928 276356
rect 112962 276308 112968 276356
rect 112874 276296 112968 276308
rect 114132 276356 114226 276368
rect 114132 276308 114138 276356
rect 114172 276308 114226 276356
rect 114132 276296 114226 276308
rect 114570 276361 114616 276373
rect 111524 276236 112624 276242
rect 111524 276202 111536 276236
rect 112612 276202 112624 276236
rect 111524 276198 112624 276202
rect 112874 276202 112922 276296
rect 114327 276291 114395 276292
rect 114570 276291 114576 276361
rect 113000 276280 114100 276286
rect 113000 276246 113012 276280
rect 114088 276246 114100 276280
rect 113000 276240 114100 276246
rect 114327 276233 114576 276291
rect 114610 276233 114616 276361
rect 114327 276231 114616 276233
rect 114327 276202 114395 276231
rect 114570 276221 114616 276231
rect 114898 276361 114944 276373
rect 114898 276233 114904 276361
rect 114938 276233 114944 276361
rect 114898 276221 114944 276233
rect 115261 276361 115307 276373
rect 115261 276233 115267 276361
rect 115301 276233 115307 276361
rect 115261 276221 115307 276233
rect 115589 276361 115635 276373
rect 115589 276233 115595 276361
rect 115629 276291 115635 276361
rect 115979 276368 116027 276458
rect 116105 276418 117205 276424
rect 116105 276384 116117 276418
rect 117193 276384 117205 276418
rect 116105 276378 117205 276384
rect 117283 276368 117331 276458
rect 115979 276356 116073 276368
rect 115979 276308 116033 276356
rect 116067 276308 116073 276356
rect 115979 276296 116073 276308
rect 117237 276356 117331 276368
rect 117237 276308 117243 276356
rect 117277 276308 117331 276356
rect 117237 276296 117331 276308
rect 115810 276291 115878 276292
rect 115629 276233 115878 276291
rect 116105 276280 117205 276286
rect 116105 276246 116117 276280
rect 117193 276246 117205 276280
rect 116105 276240 117205 276246
rect 115589 276231 115878 276233
rect 115589 276221 115635 276231
rect 112874 276198 114395 276202
rect 111524 276196 114395 276198
rect 112044 276162 114395 276196
rect 114657 276205 114857 276211
rect 114657 276171 114669 276205
rect 114845 276171 114857 276205
rect 114657 276165 114857 276171
rect 115348 276205 115548 276211
rect 115348 276171 115360 276205
rect 115536 276171 115548 276205
rect 115348 276165 115548 276171
rect 115810 276202 115878 276231
rect 117283 276202 117331 276296
rect 117461 276624 117509 276752
rect 117543 276624 117549 276752
rect 117461 276612 117549 276624
rect 118713 276752 118801 276764
rect 118713 276624 118719 276752
rect 118753 276624 118801 276752
rect 118713 276612 118801 276624
rect 120377 277105 120423 277117
rect 120377 276629 120383 277105
rect 120417 276629 120423 277105
rect 120377 276617 120423 276629
rect 120835 277105 120881 277117
rect 120835 276629 120841 277105
rect 120875 276928 120881 277105
rect 120953 277091 121018 277585
rect 121077 277413 121083 277585
rect 121117 277413 121123 277889
rect 121077 277401 121123 277413
rect 121535 277889 121605 277901
rect 121535 277413 121541 277889
rect 121575 277484 121605 277889
rect 121657 277484 121677 279396
rect 121797 279275 121849 279887
rect 122191 279275 122235 279887
rect 122360 279876 122752 279882
rect 122360 279842 122372 279876
rect 122740 279842 122752 279876
rect 122360 279836 122752 279842
rect 122808 279836 122951 279923
rect 123452 279882 123551 279923
rect 122360 279726 122951 279836
rect 122360 279720 122752 279726
rect 122360 279686 122372 279720
rect 122740 279686 122752 279720
rect 122360 279680 122752 279686
rect 122808 279639 122951 279726
rect 123060 279876 123551 279882
rect 123060 279842 123072 279876
rect 123440 279842 123551 279876
rect 123060 279720 123551 279842
rect 123060 279686 123072 279720
rect 123440 279686 123551 279720
rect 123060 279680 123551 279686
rect 123452 279639 123551 279680
rect 121797 279225 122235 279275
rect 122304 279627 122350 279639
rect 122304 279151 122310 279627
rect 122344 279151 122350 279627
rect 122304 279139 122350 279151
rect 122762 279627 123050 279639
rect 122762 279151 122768 279627
rect 122802 279151 123010 279627
rect 123044 279151 123050 279627
rect 122762 279139 123050 279151
rect 123462 279627 123551 279639
rect 123462 279151 123468 279627
rect 123502 279151 123551 279627
rect 123462 279139 123551 279151
rect 123452 279098 123551 279139
rect 122360 279092 122752 279098
rect 122360 279058 122372 279092
rect 122740 279058 122752 279092
rect 122360 279052 122752 279058
rect 123060 279092 123551 279098
rect 123060 279058 123072 279092
rect 123440 279058 123551 279092
rect 123060 279052 123551 279058
rect 122462 278353 123477 278384
rect 122418 278347 123477 278353
rect 122418 278313 122430 278347
rect 123274 278342 123477 278347
rect 123274 278313 123286 278342
rect 122418 278307 123286 278313
rect 122362 278254 122408 278266
rect 122362 277804 122368 278254
rect 122402 277804 122408 278254
rect 122362 277792 122408 277804
rect 123296 278254 123342 278266
rect 123296 277804 123302 278254
rect 123336 277804 123342 278254
rect 123296 277792 123342 277804
rect 122418 277745 123286 277751
rect 122418 277711 122430 277745
rect 123274 277711 123286 277745
rect 122418 277707 123286 277711
rect 123440 277707 123477 278342
rect 123660 278161 124206 278167
rect 123660 278127 123672 278161
rect 124194 278127 124206 278161
rect 123660 278121 124206 278127
rect 122418 277670 123477 277707
rect 121575 277413 121677 277484
rect 121535 277401 121677 277413
rect 122364 277581 123212 277587
rect 122364 277547 122432 277581
rect 123200 277547 123212 277581
rect 122364 277541 123212 277547
rect 122364 277500 122420 277541
rect 123440 277500 123477 277670
rect 123604 278068 123650 278080
rect 123604 277500 123610 278068
rect 122364 277488 122410 277500
rect 122364 277412 122370 277488
rect 122404 277412 122410 277488
rect 121133 277354 121525 277360
rect 121133 277320 121145 277354
rect 121513 277320 121525 277354
rect 121133 277198 121525 277320
rect 121133 277164 121145 277198
rect 121513 277164 121525 277198
rect 121133 277158 121525 277164
rect 121581 277117 121624 277401
rect 122364 277400 122410 277412
rect 123222 277488 123610 277500
rect 123222 277412 123228 277488
rect 123262 277412 123610 277488
rect 123222 277406 123610 277412
rect 123644 277406 123650 278068
rect 123222 277400 123650 277406
rect 122364 277359 122420 277400
rect 123604 277394 123650 277400
rect 124216 278068 124262 278080
rect 124216 277406 124222 278068
rect 124256 277528 124262 278068
rect 124256 277406 124567 277528
rect 124216 277394 124567 277406
rect 122364 277353 123212 277359
rect 122364 277319 122432 277353
rect 123200 277319 123212 277353
rect 122364 277313 123212 277319
rect 123660 277347 124206 277353
rect 123660 277313 123672 277347
rect 124194 277313 124206 277347
rect 123660 277307 124206 277313
rect 120953 276928 120958 277091
rect 120875 276809 120958 276928
rect 121013 276928 121018 277091
rect 121077 277105 121123 277117
rect 121077 276928 121083 277105
rect 121013 276809 121083 276928
rect 120875 276801 121083 276809
rect 120875 276629 120881 276801
rect 120835 276617 120881 276629
rect 121077 276629 121083 276801
rect 121117 276629 121123 277105
rect 121077 276617 121123 276629
rect 121535 277105 121624 277117
rect 121535 276629 121541 277105
rect 121575 276629 121624 277105
rect 123792 277076 123945 277307
rect 123686 277034 123945 277076
rect 123686 276881 123736 277034
rect 123913 276881 123945 277034
rect 123686 276837 123945 276881
rect 122442 276749 123828 276755
rect 122442 276715 122454 276749
rect 123816 276715 123828 276749
rect 122442 276709 123828 276715
rect 121535 276617 121624 276629
rect 122386 276656 122432 276668
rect 117461 276404 117503 276612
rect 117581 276596 118681 276602
rect 117581 276562 117593 276596
rect 118669 276562 118681 276596
rect 117581 276556 118681 276562
rect 117581 276454 118681 276460
rect 117581 276420 117593 276454
rect 118669 276420 118681 276454
rect 117581 276414 118681 276420
rect 118759 276404 118801 276612
rect 117461 276392 117549 276404
rect 117461 276264 117509 276392
rect 117543 276264 117549 276392
rect 117461 276252 117549 276264
rect 118713 276392 118801 276404
rect 118713 276264 118719 276392
rect 118753 276264 118801 276392
rect 120433 276570 120825 276576
rect 120433 276536 120445 276570
rect 120813 276536 120825 276570
rect 120433 276414 120825 276536
rect 120433 276380 120445 276414
rect 120813 276380 120825 276414
rect 120433 276374 120825 276380
rect 121133 276570 121525 276576
rect 121133 276536 121145 276570
rect 121513 276536 121525 276570
rect 121133 276414 121525 276536
rect 122386 276504 122392 276656
rect 122426 276504 122432 276656
rect 122386 276492 122432 276504
rect 123838 276656 123884 276668
rect 123838 276504 123844 276656
rect 123878 276646 123884 276656
rect 123878 276514 124112 276646
rect 123878 276504 123884 276514
rect 123838 276492 123884 276504
rect 121133 276380 121145 276414
rect 121513 276380 121525 276414
rect 122442 276445 123828 276451
rect 122442 276411 122454 276445
rect 123816 276411 123828 276445
rect 122442 276405 123828 276411
rect 121133 276374 121525 276380
rect 118713 276252 118801 276264
rect 120377 276321 120423 276333
rect 115810 276198 117331 276202
rect 117581 276236 118681 276242
rect 117581 276202 117593 276236
rect 118669 276202 118681 276236
rect 117581 276198 118681 276202
rect 115810 276196 118681 276198
rect 112719 276120 112924 276162
rect 113982 276088 114266 276098
rect 114724 276088 114783 276165
rect 113982 276085 114783 276088
rect 113982 276016 114010 276085
rect 114237 276016 114783 276085
rect 113982 275999 114783 276016
rect 115422 276088 115481 276165
rect 115810 276162 118161 276196
rect 117281 276120 117486 276162
rect 115939 276088 116223 276098
rect 115422 276085 116223 276088
rect 115422 276016 115968 276085
rect 116195 276016 116223 276085
rect 115422 275999 116223 276016
rect 113982 275998 114266 275999
rect 115939 275998 116223 275999
rect 112970 275876 114070 275882
rect 111524 275868 112624 275874
rect 111524 275834 111536 275868
rect 112612 275834 112624 275868
rect 112970 275842 112982 275876
rect 114058 275842 114070 275876
rect 116135 275876 117235 275882
rect 112970 275836 114070 275842
rect 114657 275851 114857 275857
rect 111524 275828 112624 275834
rect 111404 275806 111492 275818
rect 111404 275678 111452 275806
rect 111486 275678 111492 275806
rect 111404 275666 111492 275678
rect 112656 275806 112744 275818
rect 112656 275678 112662 275806
rect 112696 275750 112744 275806
rect 112850 275814 112938 275826
rect 112850 275750 112898 275814
rect 112696 275688 112898 275750
rect 112696 275678 112744 275688
rect 112656 275666 112744 275678
rect 111404 275458 111446 275666
rect 111524 275650 112624 275656
rect 111524 275616 111536 275650
rect 112612 275616 112624 275650
rect 111524 275610 112624 275616
rect 112702 275634 112744 275666
rect 112850 275646 112898 275688
rect 112932 275646 112938 275814
rect 112850 275634 112938 275646
rect 114102 275814 114190 275826
rect 114102 275646 114108 275814
rect 114142 275760 114190 275814
rect 114657 275817 114669 275851
rect 114845 275817 114857 275851
rect 114657 275811 114857 275817
rect 115348 275851 115548 275857
rect 115348 275817 115360 275851
rect 115536 275817 115548 275851
rect 116135 275842 116147 275876
rect 117223 275842 117235 275876
rect 116135 275836 117235 275842
rect 117581 275868 118681 275874
rect 117581 275834 117593 275868
rect 118669 275834 118681 275868
rect 117581 275828 118681 275834
rect 120377 275845 120383 276321
rect 120417 275845 120423 276321
rect 120377 275833 120423 275845
rect 120835 276321 120881 276333
rect 120835 275845 120841 276321
rect 120875 276139 120881 276321
rect 121077 276321 121123 276333
rect 121077 276139 121083 276321
rect 120875 276118 121083 276139
rect 120875 276054 120958 276118
rect 121014 276054 121083 276118
rect 120875 276032 121083 276054
rect 120875 275845 120881 276032
rect 120835 275833 120881 275845
rect 115348 275811 115548 275817
rect 116015 275814 116103 275826
rect 114570 275789 114616 275801
rect 114570 275760 114576 275789
rect 114142 275646 114576 275760
rect 114102 275634 114576 275646
rect 111524 275508 112624 275514
rect 111524 275474 111536 275508
rect 112612 275474 112624 275508
rect 111524 275468 112624 275474
rect 112702 275458 112746 275634
rect 111404 275446 111492 275458
rect 111404 275318 111452 275446
rect 111486 275318 111492 275446
rect 111404 275306 111492 275318
rect 112656 275446 112746 275458
rect 112656 275318 112662 275446
rect 112696 275414 112746 275446
rect 112850 275534 112892 275634
rect 114148 275627 114576 275634
rect 112970 275618 114070 275624
rect 112970 275584 112982 275618
rect 114058 275584 114070 275618
rect 112970 275578 114070 275584
rect 114148 275534 114190 275627
rect 112850 275496 114190 275534
rect 112696 275366 112744 275414
rect 112850 275402 112892 275496
rect 112970 275452 114070 275458
rect 112970 275418 112982 275452
rect 114058 275418 114070 275452
rect 112970 275412 114070 275418
rect 114148 275402 114190 275496
rect 114570 275421 114576 275627
rect 114610 275421 114616 275789
rect 114570 275409 114616 275421
rect 114898 275789 114944 275801
rect 114898 275421 114904 275789
rect 114938 275421 114944 275789
rect 114898 275409 114944 275421
rect 115261 275789 115307 275801
rect 115261 275421 115267 275789
rect 115301 275421 115307 275789
rect 115261 275409 115307 275421
rect 115589 275789 115635 275801
rect 115589 275421 115595 275789
rect 115629 275760 115635 275789
rect 116015 275760 116063 275814
rect 115629 275646 116063 275760
rect 116097 275646 116103 275814
rect 115629 275634 116103 275646
rect 117267 275814 117355 275826
rect 117267 275646 117273 275814
rect 117307 275750 117355 275814
rect 117461 275806 117549 275818
rect 117461 275750 117509 275806
rect 117307 275688 117509 275750
rect 117307 275646 117355 275688
rect 117267 275634 117355 275646
rect 117461 275678 117509 275688
rect 117543 275678 117549 275806
rect 117461 275666 117549 275678
rect 118713 275806 118801 275818
rect 118713 275678 118719 275806
rect 118753 275678 118801 275806
rect 118713 275666 118801 275678
rect 117461 275634 117503 275666
rect 115629 275627 116057 275634
rect 115629 275421 115635 275627
rect 115589 275409 115635 275421
rect 116015 275534 116057 275627
rect 116135 275618 117235 275624
rect 116135 275584 116147 275618
rect 117223 275584 117235 275618
rect 116135 275578 117235 275584
rect 117313 275534 117355 275634
rect 116015 275496 117355 275534
rect 112850 275390 112938 275402
rect 112850 275366 112898 275390
rect 112696 275318 112898 275366
rect 112656 275306 112898 275318
rect 111404 275098 111446 275306
rect 112702 275304 112898 275306
rect 111524 275290 112624 275296
rect 111524 275256 111536 275290
rect 112612 275256 112624 275290
rect 111524 275250 112624 275256
rect 111524 275148 112624 275154
rect 111524 275114 111536 275148
rect 112612 275114 112624 275148
rect 111524 275108 112624 275114
rect 112702 275098 112744 275304
rect 112850 275222 112898 275304
rect 112932 275222 112938 275390
rect 112850 275210 112938 275222
rect 114102 275390 114190 275402
rect 116015 275402 116057 275496
rect 116135 275452 117235 275458
rect 116135 275418 116147 275452
rect 117223 275418 117235 275452
rect 116135 275412 117235 275418
rect 117313 275402 117355 275496
rect 117459 275458 117503 275634
rect 117581 275650 118681 275656
rect 117581 275616 117593 275650
rect 118669 275616 118681 275650
rect 117581 275610 118681 275616
rect 117581 275508 118681 275514
rect 117581 275474 117593 275508
rect 118669 275474 118681 275508
rect 117581 275468 118681 275474
rect 118759 275458 118801 275666
rect 120433 275786 120825 275792
rect 120433 275752 120445 275786
rect 120813 275752 120825 275786
rect 120433 275630 120825 275752
rect 120433 275596 120445 275630
rect 120813 275596 120825 275630
rect 120433 275590 120825 275596
rect 117459 275446 117549 275458
rect 117459 275414 117509 275446
rect 114102 275222 114108 275390
rect 114142 275222 114190 275390
rect 114657 275393 114857 275399
rect 114657 275359 114669 275393
rect 114845 275359 114857 275393
rect 114657 275353 114857 275359
rect 115348 275393 115548 275399
rect 115348 275359 115360 275393
rect 115536 275359 115548 275393
rect 115348 275353 115548 275359
rect 116015 275390 116103 275402
rect 114720 275285 114790 275353
rect 114102 275210 114190 275222
rect 114308 275201 114790 275285
rect 114865 275296 114970 275313
rect 114865 275228 114885 275296
rect 114948 275228 114970 275296
rect 114865 275206 114970 275228
rect 115235 275296 115340 275313
rect 115235 275228 115257 275296
rect 115320 275228 115340 275296
rect 115235 275206 115340 275228
rect 115415 275285 115485 275353
rect 112970 275194 114070 275200
rect 112970 275160 112982 275194
rect 114058 275160 114070 275194
rect 112970 275154 114070 275160
rect 111404 275086 111492 275098
rect 111404 274958 111452 275086
rect 111486 274958 111492 275086
rect 111404 274946 111492 274958
rect 112656 275086 112744 275098
rect 114308 275086 114343 275201
rect 114720 275171 114790 275201
rect 115415 275201 115897 275285
rect 116015 275222 116063 275390
rect 116097 275222 116103 275390
rect 116015 275210 116103 275222
rect 117267 275390 117355 275402
rect 117267 275222 117273 275390
rect 117307 275366 117355 275390
rect 117461 275366 117509 275414
rect 117307 275318 117509 275366
rect 117543 275318 117549 275446
rect 117307 275306 117549 275318
rect 118713 275446 118801 275458
rect 118713 275318 118719 275446
rect 118753 275318 118801 275446
rect 118713 275306 118801 275318
rect 117307 275304 117503 275306
rect 117307 275222 117355 275304
rect 117267 275210 117355 275222
rect 115415 275171 115485 275201
rect 114657 275165 114857 275171
rect 114657 275131 114669 275165
rect 114845 275131 114857 275165
rect 114657 275125 114857 275131
rect 115348 275165 115548 275171
rect 115348 275131 115360 275165
rect 115536 275131 115548 275165
rect 115348 275125 115548 275131
rect 112656 274958 112662 275086
rect 112696 274958 112744 275086
rect 113843 275056 114343 275086
rect 113000 275050 114343 275056
rect 113000 275016 113012 275050
rect 114088 275045 114343 275050
rect 114570 275103 114616 275115
rect 114088 275016 114100 275045
rect 113000 275010 114100 275016
rect 112656 274946 112744 274958
rect 111404 274738 111446 274946
rect 111524 274930 112624 274936
rect 111524 274896 111536 274930
rect 112612 274896 112624 274930
rect 111524 274890 112624 274896
rect 111524 274788 112624 274794
rect 111524 274754 111536 274788
rect 112612 274754 112624 274788
rect 111524 274748 112624 274754
rect 112702 274738 112744 274946
rect 111404 274726 111492 274738
rect 111404 274598 111452 274726
rect 111486 274598 111492 274726
rect 111404 274586 111492 274598
rect 112656 274726 112744 274738
rect 112656 274598 112662 274726
rect 112696 274598 112744 274726
rect 112656 274586 112744 274598
rect 112874 274988 112968 275000
rect 112874 274940 112928 274988
rect 112962 274940 112968 274988
rect 112874 274928 112968 274940
rect 114132 274988 114226 275000
rect 114132 274940 114138 274988
rect 114172 274940 114226 274988
rect 114132 274928 114226 274940
rect 112874 274836 112922 274928
rect 113000 274912 114100 274918
rect 113000 274878 113012 274912
rect 114088 274878 114100 274912
rect 113000 274872 114100 274878
rect 114178 274836 114226 274928
rect 112874 274792 114226 274836
rect 114324 274978 114396 274994
rect 114324 274895 114342 274978
rect 114377 274895 114396 274978
rect 114570 274975 114576 275103
rect 114610 274975 114616 275103
rect 114570 274963 114616 274975
rect 114898 275103 114944 275115
rect 114898 274975 114904 275103
rect 114938 274975 114944 275103
rect 114898 274963 114944 274975
rect 115261 275103 115307 275115
rect 115261 274975 115267 275103
rect 115301 274975 115307 275103
rect 115261 274963 115307 274975
rect 115589 275103 115635 275115
rect 115589 274975 115595 275103
rect 115629 274975 115635 275103
rect 115862 275086 115897 275201
rect 116135 275194 117235 275200
rect 116135 275160 116147 275194
rect 117223 275160 117235 275194
rect 116135 275154 117235 275160
rect 117461 275098 117503 275304
rect 117581 275290 118681 275296
rect 117581 275256 117593 275290
rect 118669 275256 118681 275290
rect 117581 275250 118681 275256
rect 117581 275148 118681 275154
rect 117581 275114 117593 275148
rect 118669 275114 118681 275148
rect 117581 275108 118681 275114
rect 118759 275098 118801 275306
rect 117461 275086 117549 275098
rect 115862 275056 116362 275086
rect 115862 275050 117205 275056
rect 115862 275045 116117 275050
rect 116105 275016 116117 275045
rect 117193 275016 117205 275050
rect 116105 275010 117205 275016
rect 115589 274963 115635 274975
rect 115809 274978 115881 274994
rect 114657 274947 114857 274953
rect 114657 274913 114669 274947
rect 114845 274913 114857 274947
rect 114657 274907 114857 274913
rect 115348 274947 115548 274953
rect 115348 274913 115360 274947
rect 115536 274913 115548 274947
rect 115348 274907 115548 274913
rect 114324 274863 114396 274895
rect 115809 274895 115828 274978
rect 115863 274895 115881 274978
rect 114843 274863 115030 274878
rect 114324 274818 114781 274863
rect 112874 274702 112922 274792
rect 113000 274752 114100 274758
rect 113000 274718 113012 274752
rect 114088 274718 114100 274752
rect 113000 274712 114100 274718
rect 114178 274702 114226 274792
rect 114737 274763 114781 274818
rect 114843 274811 114868 274863
rect 114966 274811 115030 274863
rect 114843 274793 115030 274811
rect 115175 274863 115362 274878
rect 115809 274863 115881 274895
rect 115175 274811 115239 274863
rect 115337 274811 115362 274863
rect 115175 274793 115362 274811
rect 115424 274818 115881 274863
rect 115979 274988 116073 275000
rect 115979 274940 116033 274988
rect 116067 274940 116073 274988
rect 115979 274928 116073 274940
rect 117237 274988 117331 275000
rect 117237 274940 117243 274988
rect 117277 274940 117331 274988
rect 117237 274928 117331 274940
rect 115979 274836 116027 274928
rect 116105 274912 117205 274918
rect 116105 274878 116117 274912
rect 117193 274878 117205 274912
rect 116105 274872 117205 274878
rect 117283 274836 117331 274928
rect 115424 274763 115468 274818
rect 115979 274792 117331 274836
rect 114657 274757 114857 274763
rect 114657 274723 114669 274757
rect 114845 274723 114857 274757
rect 114657 274717 114857 274723
rect 115348 274757 115548 274763
rect 115348 274723 115360 274757
rect 115536 274723 115548 274757
rect 115348 274717 115548 274723
rect 112874 274690 112968 274702
rect 112874 274642 112928 274690
rect 112962 274642 112968 274690
rect 112874 274630 112968 274642
rect 114132 274690 114226 274702
rect 114132 274642 114138 274690
rect 114172 274642 114226 274690
rect 114132 274630 114226 274642
rect 114570 274695 114616 274707
rect 111524 274570 112624 274576
rect 111524 274536 111536 274570
rect 112612 274536 112624 274570
rect 111524 274532 112624 274536
rect 112874 274536 112922 274630
rect 114327 274625 114395 274626
rect 114570 274625 114576 274695
rect 113000 274614 114100 274620
rect 113000 274580 113012 274614
rect 114088 274580 114100 274614
rect 113000 274574 114100 274580
rect 114327 274567 114576 274625
rect 114610 274567 114616 274695
rect 114327 274565 114616 274567
rect 114327 274536 114395 274565
rect 114570 274555 114616 274565
rect 114898 274695 114944 274707
rect 114898 274567 114904 274695
rect 114938 274567 114944 274695
rect 114898 274555 114944 274567
rect 115261 274695 115307 274707
rect 115261 274567 115267 274695
rect 115301 274567 115307 274695
rect 115261 274555 115307 274567
rect 115589 274695 115635 274707
rect 115589 274567 115595 274695
rect 115629 274625 115635 274695
rect 115979 274702 116027 274792
rect 116105 274752 117205 274758
rect 116105 274718 116117 274752
rect 117193 274718 117205 274752
rect 116105 274712 117205 274718
rect 117283 274702 117331 274792
rect 115979 274690 116073 274702
rect 115979 274642 116033 274690
rect 116067 274642 116073 274690
rect 115979 274630 116073 274642
rect 117237 274690 117331 274702
rect 117237 274642 117243 274690
rect 117277 274642 117331 274690
rect 117237 274630 117331 274642
rect 115810 274625 115878 274626
rect 115629 274567 115878 274625
rect 116105 274614 117205 274620
rect 116105 274580 116117 274614
rect 117193 274580 117205 274614
rect 116105 274574 117205 274580
rect 115589 274565 115878 274567
rect 115589 274555 115635 274565
rect 112874 274532 114395 274536
rect 111524 274530 114395 274532
rect 108355 274505 111012 274509
rect 106072 274503 111014 274505
rect 102557 274070 105283 274145
rect 102557 273772 102621 274070
rect 105204 273772 105283 274070
rect 106053 274267 111014 274503
rect 112044 274496 114395 274530
rect 114657 274539 114857 274545
rect 114657 274505 114669 274539
rect 114845 274505 114857 274539
rect 114657 274499 114857 274505
rect 115348 274539 115548 274545
rect 115348 274505 115360 274539
rect 115536 274505 115548 274539
rect 115348 274499 115548 274505
rect 115810 274536 115878 274565
rect 117283 274536 117331 274630
rect 117461 274958 117509 275086
rect 117543 274958 117549 275086
rect 117461 274946 117549 274958
rect 118713 275086 118801 275098
rect 118713 274958 118719 275086
rect 118753 274958 118801 275086
rect 120377 275537 120423 275549
rect 120377 275061 120383 275537
rect 120417 275061 120423 275537
rect 120377 275049 120423 275061
rect 120835 275537 120881 275549
rect 120835 275061 120841 275537
rect 120875 275061 120881 275537
rect 120835 275049 120881 275061
rect 118713 274946 118801 274958
rect 117461 274738 117503 274946
rect 117581 274930 118681 274936
rect 117581 274896 117593 274930
rect 118669 274896 118681 274930
rect 117581 274890 118681 274896
rect 117581 274788 118681 274794
rect 117581 274754 117593 274788
rect 118669 274754 118681 274788
rect 117581 274748 118681 274754
rect 118759 274738 118801 274946
rect 120433 275002 120825 275008
rect 120433 274968 120445 275002
rect 120813 274968 120825 275002
rect 120433 274846 120825 274968
rect 120433 274812 120445 274846
rect 120813 274812 120825 274846
rect 120433 274806 120825 274812
rect 117461 274726 117549 274738
rect 117461 274598 117509 274726
rect 117543 274598 117549 274726
rect 117461 274586 117549 274598
rect 118713 274726 118801 274738
rect 118713 274598 118719 274726
rect 118753 274598 118801 274726
rect 118713 274586 118801 274598
rect 120377 274753 120423 274765
rect 115810 274532 117331 274536
rect 117581 274570 118681 274576
rect 117581 274536 117593 274570
rect 118669 274536 118681 274570
rect 117581 274532 118681 274536
rect 115810 274530 118681 274532
rect 112719 274454 112924 274496
rect 113982 274422 114266 274432
rect 114724 274422 114783 274499
rect 113982 274419 114783 274422
rect 113982 274350 114010 274419
rect 114237 274350 114783 274419
rect 113982 274333 114783 274350
rect 115422 274422 115481 274499
rect 115810 274496 118161 274530
rect 117281 274454 117486 274496
rect 115939 274422 116223 274432
rect 115422 274419 116223 274422
rect 115422 274350 115968 274419
rect 116195 274350 116223 274419
rect 115422 274333 116223 274350
rect 113982 274332 114266 274333
rect 115939 274332 116223 274333
rect 120377 274277 120383 274753
rect 120417 274277 120423 274753
rect 106053 273841 111015 274267
rect 120377 274265 120423 274277
rect 120835 274753 120881 274765
rect 120835 274277 120841 274753
rect 120875 274277 120881 274753
rect 120835 274265 120881 274277
rect 120433 274218 120825 274224
rect 112970 274210 114070 274216
rect 111524 274202 112624 274208
rect 111524 274168 111536 274202
rect 112612 274168 112624 274202
rect 112970 274176 112982 274210
rect 114058 274176 114070 274210
rect 116135 274210 117235 274216
rect 112970 274170 114070 274176
rect 114657 274185 114857 274191
rect 111524 274162 112624 274168
rect 111404 274140 111492 274152
rect 111404 274012 111452 274140
rect 111486 274012 111492 274140
rect 111404 274000 111492 274012
rect 112656 274140 112744 274152
rect 112656 274012 112662 274140
rect 112696 274084 112744 274140
rect 112850 274148 112938 274160
rect 112850 274084 112898 274148
rect 112696 274022 112898 274084
rect 112696 274012 112744 274022
rect 112656 274000 112744 274012
rect 102557 273716 105283 273772
rect 108199 273428 108478 273841
rect 105964 273149 108478 273428
rect 111404 273792 111446 274000
rect 111524 273984 112624 273990
rect 111524 273950 111536 273984
rect 112612 273950 112624 273984
rect 111524 273944 112624 273950
rect 112702 273968 112744 274000
rect 112850 273980 112898 274022
rect 112932 273980 112938 274148
rect 112850 273968 112938 273980
rect 114102 274148 114190 274160
rect 114102 273980 114108 274148
rect 114142 274094 114190 274148
rect 114657 274151 114669 274185
rect 114845 274151 114857 274185
rect 114657 274145 114857 274151
rect 115348 274185 115548 274191
rect 115348 274151 115360 274185
rect 115536 274151 115548 274185
rect 116135 274176 116147 274210
rect 117223 274176 117235 274210
rect 116135 274170 117235 274176
rect 117581 274202 118681 274208
rect 117581 274168 117593 274202
rect 118669 274168 118681 274202
rect 117581 274162 118681 274168
rect 120433 274184 120445 274218
rect 120813 274184 120825 274218
rect 115348 274145 115548 274151
rect 116015 274148 116103 274160
rect 114570 274123 114616 274135
rect 114570 274094 114576 274123
rect 114142 273980 114576 274094
rect 114102 273968 114576 273980
rect 111524 273842 112624 273848
rect 111524 273808 111536 273842
rect 112612 273808 112624 273842
rect 111524 273802 112624 273808
rect 112702 273792 112746 273968
rect 111404 273780 111492 273792
rect 111404 273652 111452 273780
rect 111486 273652 111492 273780
rect 111404 273640 111492 273652
rect 112656 273780 112746 273792
rect 112656 273652 112662 273780
rect 112696 273748 112746 273780
rect 112850 273868 112892 273968
rect 114148 273961 114576 273968
rect 112970 273952 114070 273958
rect 112970 273918 112982 273952
rect 114058 273918 114070 273952
rect 112970 273912 114070 273918
rect 114148 273868 114190 273961
rect 112850 273830 114190 273868
rect 112696 273700 112744 273748
rect 112850 273736 112892 273830
rect 112970 273786 114070 273792
rect 112970 273752 112982 273786
rect 114058 273752 114070 273786
rect 112970 273746 114070 273752
rect 114148 273736 114190 273830
rect 114570 273755 114576 273961
rect 114610 273755 114616 274123
rect 114570 273743 114616 273755
rect 114898 274123 114944 274135
rect 114898 273755 114904 274123
rect 114938 273755 114944 274123
rect 114898 273743 114944 273755
rect 115261 274123 115307 274135
rect 115261 273755 115267 274123
rect 115301 273755 115307 274123
rect 115261 273743 115307 273755
rect 115589 274123 115635 274135
rect 115589 273755 115595 274123
rect 115629 274094 115635 274123
rect 116015 274094 116063 274148
rect 115629 273980 116063 274094
rect 116097 273980 116103 274148
rect 115629 273968 116103 273980
rect 117267 274148 117355 274160
rect 117267 273980 117273 274148
rect 117307 274084 117355 274148
rect 117461 274140 117549 274152
rect 117461 274084 117509 274140
rect 117307 274022 117509 274084
rect 117307 273980 117355 274022
rect 117267 273968 117355 273980
rect 117461 274012 117509 274022
rect 117543 274012 117549 274140
rect 117461 274000 117549 274012
rect 118713 274140 118801 274152
rect 118713 274012 118719 274140
rect 118753 274012 118801 274140
rect 120433 274062 120825 274184
rect 120433 274028 120445 274062
rect 120813 274028 120825 274062
rect 120433 274022 120825 274028
rect 118713 274000 118801 274012
rect 117461 273968 117503 274000
rect 115629 273961 116057 273968
rect 115629 273755 115635 273961
rect 115589 273743 115635 273755
rect 116015 273868 116057 273961
rect 116135 273952 117235 273958
rect 116135 273918 116147 273952
rect 117223 273918 117235 273952
rect 116135 273912 117235 273918
rect 117313 273868 117355 273968
rect 116015 273830 117355 273868
rect 112850 273724 112938 273736
rect 112850 273700 112898 273724
rect 112696 273652 112898 273700
rect 112656 273640 112898 273652
rect 111404 273432 111446 273640
rect 112702 273638 112898 273640
rect 111524 273624 112624 273630
rect 111524 273590 111536 273624
rect 112612 273590 112624 273624
rect 111524 273584 112624 273590
rect 111524 273482 112624 273488
rect 111524 273448 111536 273482
rect 112612 273448 112624 273482
rect 111524 273442 112624 273448
rect 112702 273432 112744 273638
rect 112850 273556 112898 273638
rect 112932 273556 112938 273724
rect 112850 273544 112938 273556
rect 114102 273724 114190 273736
rect 116015 273736 116057 273830
rect 116135 273786 117235 273792
rect 116135 273752 116147 273786
rect 117223 273752 117235 273786
rect 116135 273746 117235 273752
rect 117313 273736 117355 273830
rect 117459 273792 117503 273968
rect 117581 273984 118681 273990
rect 117581 273950 117593 273984
rect 118669 273950 118681 273984
rect 117581 273944 118681 273950
rect 117581 273842 118681 273848
rect 117581 273808 117593 273842
rect 118669 273808 118681 273842
rect 117581 273802 118681 273808
rect 118759 273792 118801 274000
rect 117459 273780 117549 273792
rect 117459 273748 117509 273780
rect 114102 273556 114108 273724
rect 114142 273556 114190 273724
rect 114657 273727 114857 273733
rect 114657 273693 114669 273727
rect 114845 273693 114857 273727
rect 114657 273687 114857 273693
rect 115348 273727 115548 273733
rect 115348 273693 115360 273727
rect 115536 273693 115548 273727
rect 115348 273687 115548 273693
rect 116015 273724 116103 273736
rect 114720 273619 114790 273687
rect 114102 273544 114190 273556
rect 114308 273535 114790 273619
rect 114865 273630 114970 273647
rect 114865 273562 114885 273630
rect 114948 273562 114970 273630
rect 114865 273540 114970 273562
rect 115235 273630 115340 273647
rect 115235 273562 115257 273630
rect 115320 273562 115340 273630
rect 115235 273540 115340 273562
rect 115415 273619 115485 273687
rect 112970 273528 114070 273534
rect 112970 273494 112982 273528
rect 114058 273494 114070 273528
rect 112970 273488 114070 273494
rect 111404 273420 111492 273432
rect 111404 273292 111452 273420
rect 111486 273292 111492 273420
rect 111404 273280 111492 273292
rect 112656 273420 112744 273432
rect 114308 273420 114343 273535
rect 114720 273505 114790 273535
rect 115415 273535 115897 273619
rect 116015 273556 116063 273724
rect 116097 273556 116103 273724
rect 116015 273544 116103 273556
rect 117267 273724 117355 273736
rect 117267 273556 117273 273724
rect 117307 273700 117355 273724
rect 117461 273700 117509 273748
rect 117307 273652 117509 273700
rect 117543 273652 117549 273780
rect 117307 273640 117549 273652
rect 118713 273780 118801 273792
rect 118713 273652 118719 273780
rect 118753 273652 118801 273780
rect 118713 273640 118801 273652
rect 117307 273638 117503 273640
rect 117307 273556 117355 273638
rect 117267 273544 117355 273556
rect 115415 273505 115485 273535
rect 114657 273499 114857 273505
rect 114657 273465 114669 273499
rect 114845 273465 114857 273499
rect 114657 273459 114857 273465
rect 115348 273499 115548 273505
rect 115348 273465 115360 273499
rect 115536 273465 115548 273499
rect 115348 273459 115548 273465
rect 112656 273292 112662 273420
rect 112696 273292 112744 273420
rect 113843 273390 114343 273420
rect 113000 273384 114343 273390
rect 113000 273350 113012 273384
rect 114088 273379 114343 273384
rect 114570 273437 114616 273449
rect 114088 273350 114100 273379
rect 113000 273344 114100 273350
rect 112656 273280 112744 273292
rect 105964 270099 106243 273149
rect 111404 273072 111446 273280
rect 111524 273264 112624 273270
rect 111524 273230 111536 273264
rect 112612 273230 112624 273264
rect 111524 273224 112624 273230
rect 111524 273122 112624 273128
rect 111524 273088 111536 273122
rect 112612 273088 112624 273122
rect 111524 273082 112624 273088
rect 112702 273072 112744 273280
rect 111404 273060 111492 273072
rect 111404 272932 111452 273060
rect 111486 272932 111492 273060
rect 111404 272920 111492 272932
rect 112656 273060 112744 273072
rect 112656 272932 112662 273060
rect 112696 272932 112744 273060
rect 112656 272920 112744 272932
rect 112874 273322 112968 273334
rect 112874 273274 112928 273322
rect 112962 273274 112968 273322
rect 112874 273262 112968 273274
rect 114132 273322 114226 273334
rect 114132 273274 114138 273322
rect 114172 273274 114226 273322
rect 114132 273262 114226 273274
rect 112874 273170 112922 273262
rect 113000 273246 114100 273252
rect 113000 273212 113012 273246
rect 114088 273212 114100 273246
rect 113000 273206 114100 273212
rect 114178 273170 114226 273262
rect 112874 273126 114226 273170
rect 114324 273312 114396 273328
rect 114324 273229 114342 273312
rect 114377 273229 114396 273312
rect 114570 273309 114576 273437
rect 114610 273309 114616 273437
rect 114570 273297 114616 273309
rect 114898 273437 114944 273449
rect 114898 273309 114904 273437
rect 114938 273309 114944 273437
rect 114898 273297 114944 273309
rect 115261 273437 115307 273449
rect 115261 273309 115267 273437
rect 115301 273309 115307 273437
rect 115261 273297 115307 273309
rect 115589 273437 115635 273449
rect 115589 273309 115595 273437
rect 115629 273309 115635 273437
rect 115862 273420 115897 273535
rect 116135 273528 117235 273534
rect 116135 273494 116147 273528
rect 117223 273494 117235 273528
rect 116135 273488 117235 273494
rect 117461 273432 117503 273638
rect 117581 273624 118681 273630
rect 117581 273590 117593 273624
rect 118669 273590 118681 273624
rect 117581 273584 118681 273590
rect 117581 273482 118681 273488
rect 117581 273448 117593 273482
rect 118669 273448 118681 273482
rect 117581 273442 118681 273448
rect 118759 273432 118801 273640
rect 120377 273969 120423 273981
rect 120377 273493 120383 273969
rect 120417 273493 120423 273969
rect 120377 273481 120423 273493
rect 120835 273969 120881 273981
rect 120835 273493 120841 273969
rect 120875 273778 120881 273969
rect 120950 273778 121028 276032
rect 121077 275845 121083 276032
rect 121117 275845 121123 276321
rect 121077 275833 121123 275845
rect 121535 276321 121581 276333
rect 121535 275845 121541 276321
rect 121575 276135 121581 276321
rect 121802 276227 121933 276287
rect 121802 276172 121822 276227
rect 121801 276135 121822 276172
rect 121575 276028 121822 276135
rect 121575 275845 121581 276028
rect 121802 276007 121822 276028
rect 121912 276007 121933 276227
rect 122096 276131 122427 276154
rect 122096 276060 122120 276131
rect 122404 276118 122427 276131
rect 124055 276118 124112 276514
rect 122404 276060 124349 276118
rect 122096 276049 124349 276060
rect 124445 276083 124567 277394
rect 122096 276035 122427 276049
rect 121802 275945 121933 276007
rect 121535 275833 121581 275845
rect 122390 275807 122422 276035
rect 122629 275863 122686 276049
rect 122466 275857 122866 275863
rect 122466 275823 122478 275857
rect 122854 275823 122866 275857
rect 122466 275817 122866 275823
rect 122970 275807 123002 276049
rect 123272 275863 123329 276049
rect 123102 275857 123502 275863
rect 123102 275823 123114 275857
rect 123490 275823 123502 275857
rect 123102 275817 123502 275823
rect 123605 275807 123637 276049
rect 123915 275863 123972 276049
rect 124240 275863 124272 276049
rect 124445 275982 124465 276083
rect 124549 275982 124567 276083
rect 124445 275955 124567 275982
rect 123738 275857 124138 275863
rect 123738 275823 123750 275857
rect 124126 275823 124138 275857
rect 123738 275817 124138 275823
rect 124240 275857 124774 275863
rect 124240 275823 124386 275857
rect 124762 275823 124774 275857
rect 124240 275817 124774 275823
rect 124240 275807 124374 275817
rect 122379 275795 122425 275807
rect 121133 275786 121525 275792
rect 121133 275752 121145 275786
rect 121513 275752 121525 275786
rect 121133 275630 121525 275752
rect 122379 275727 122385 275795
rect 122419 275727 122425 275795
rect 122379 275715 122425 275727
rect 122907 275795 123061 275807
rect 122907 275727 122913 275795
rect 122947 275727 123021 275795
rect 123055 275727 123061 275795
rect 122907 275715 123061 275727
rect 123543 275795 123697 275807
rect 123543 275727 123549 275795
rect 123583 275727 123657 275795
rect 123691 275727 123697 275795
rect 123543 275715 123697 275727
rect 124179 275797 124374 275807
rect 124179 275795 124333 275797
rect 124179 275727 124185 275795
rect 124219 275727 124293 275795
rect 124327 275727 124333 275795
rect 124179 275715 124333 275727
rect 124815 275795 124861 275807
rect 124815 275727 124821 275795
rect 124855 275727 124861 275795
rect 124815 275715 124861 275727
rect 122466 275699 122866 275705
rect 122466 275665 122478 275699
rect 122854 275665 122866 275699
rect 122466 275659 122866 275665
rect 123102 275699 123502 275705
rect 123102 275665 123114 275699
rect 123490 275665 123502 275699
rect 123102 275659 123502 275665
rect 123738 275699 124138 275705
rect 123738 275665 123750 275699
rect 124126 275665 124138 275699
rect 123738 275659 124138 275665
rect 121133 275596 121145 275630
rect 121513 275596 121525 275630
rect 121133 275590 121525 275596
rect 121077 275537 121123 275549
rect 121077 275061 121083 275537
rect 121117 275061 121123 275537
rect 121077 275049 121123 275061
rect 121535 275537 121628 275549
rect 121535 275061 121541 275537
rect 121575 275070 121628 275537
rect 124244 275475 124285 275715
rect 124374 275699 124774 275705
rect 124374 275665 124386 275699
rect 124762 275665 124774 275699
rect 124374 275659 124774 275665
rect 124818 275475 124859 275715
rect 124244 275432 124859 275475
rect 123213 275386 123457 275431
rect 122354 275289 122587 275333
rect 122354 275070 122391 275289
rect 121575 275061 122391 275070
rect 121535 275049 122391 275061
rect 121133 275002 121525 275008
rect 121133 274968 121145 275002
rect 121513 274968 121525 275002
rect 121133 274846 121525 274968
rect 121133 274812 121145 274846
rect 121513 274812 121525 274846
rect 121133 274806 121525 274812
rect 121581 274783 122391 275049
rect 122556 274783 122587 275289
rect 123213 275173 123245 275386
rect 123426 275336 123457 275386
rect 123426 275231 124318 275336
rect 123426 275173 123457 275231
rect 123213 275140 123457 275173
rect 124132 274973 124318 275231
rect 123881 274943 124318 274973
rect 125452 275158 128452 275523
rect 123881 274940 124366 274943
rect 122956 274934 123948 274940
rect 122956 274900 122968 274934
rect 123936 274900 123948 274934
rect 122956 274894 123948 274900
rect 122900 274850 122946 274862
rect 122900 274807 122906 274850
rect 121581 274765 122587 274783
rect 121077 274753 121123 274765
rect 121077 274277 121083 274753
rect 121117 274277 121123 274753
rect 121077 274265 121123 274277
rect 121535 274753 122587 274765
rect 121535 274277 121541 274753
rect 121575 274736 122587 274753
rect 122706 274765 122906 274807
rect 121575 274277 121628 274736
rect 122706 274454 122746 274765
rect 122900 274674 122906 274765
rect 122940 274674 122946 274850
rect 122900 274662 122946 274674
rect 123958 274850 124004 274862
rect 123958 274674 123964 274850
rect 123998 274674 124004 274850
rect 123958 274662 124004 274674
rect 122956 274624 123948 274630
rect 122956 274590 122968 274624
rect 123936 274590 123948 274624
rect 122956 274584 123948 274590
rect 124116 274584 124366 274940
rect 123879 274574 124366 274584
rect 123879 274551 124148 274574
rect 122706 274452 123624 274454
rect 122706 274445 123670 274452
rect 122706 274418 123527 274445
rect 123497 274408 123527 274418
rect 123647 274408 123670 274445
rect 123497 274401 123670 274408
rect 124001 274397 124921 274447
rect 124001 274356 124100 274397
rect 122281 274350 122477 274356
rect 122281 274316 122293 274350
rect 122461 274316 122477 274350
rect 122281 274310 122477 274316
rect 122697 274350 124137 274356
rect 122697 274316 122709 274350
rect 122877 274316 123125 274350
rect 123293 274316 123541 274350
rect 123709 274316 123957 274350
rect 124125 274316 124137 274350
rect 122697 274310 124137 274316
rect 124357 274350 124553 274356
rect 124357 274316 124373 274350
rect 124541 274316 124553 274350
rect 124357 274310 124553 274316
rect 121535 274265 121628 274277
rect 122225 274266 122271 274278
rect 121133 274218 121525 274224
rect 121133 274184 121145 274218
rect 121513 274184 121525 274218
rect 121133 274062 121525 274184
rect 121133 274028 121145 274062
rect 121513 274028 121525 274062
rect 121133 274022 121525 274028
rect 121077 273969 121123 273981
rect 121077 273778 121083 273969
rect 120875 273756 121083 273778
rect 120875 273692 120961 273756
rect 121017 273692 121083 273756
rect 120875 273671 121083 273692
rect 120875 273493 120881 273671
rect 120835 273481 120881 273493
rect 121077 273493 121083 273671
rect 121117 273493 121123 273969
rect 121077 273481 121123 273493
rect 121535 273969 121581 273981
rect 121535 273493 121541 273969
rect 121575 273769 121581 273969
rect 121803 273825 121934 273885
rect 121803 273770 121823 273825
rect 121764 273769 121823 273770
rect 121575 273662 121823 273769
rect 121575 273493 121581 273662
rect 121764 273661 121823 273662
rect 121803 273605 121823 273661
rect 121913 273605 121934 273825
rect 122225 273790 122231 274266
rect 122265 273790 122271 274266
rect 122225 273778 122271 273790
rect 122483 274266 122529 274278
rect 122483 273790 122489 274266
rect 122523 273790 122529 274266
rect 122641 274266 122687 274278
rect 122641 274044 122647 274266
rect 122483 273778 122529 273790
rect 122602 273790 122647 274044
rect 122681 273790 122687 274266
rect 122602 273778 122687 273790
rect 122899 274266 122945 274278
rect 122899 273790 122905 274266
rect 122939 273790 122945 274266
rect 123057 274266 123103 274278
rect 123057 274044 123063 274266
rect 122899 273778 122945 273790
rect 123018 273790 123063 274044
rect 123097 273790 123103 274266
rect 123018 273778 123103 273790
rect 123315 274266 123361 274278
rect 123315 273790 123321 274266
rect 123355 273790 123361 274266
rect 123473 274266 123519 274278
rect 123473 274044 123479 274266
rect 123315 273778 123361 273790
rect 123434 273790 123479 274044
rect 123513 273790 123519 274266
rect 123434 273778 123519 273790
rect 123731 274266 123777 274278
rect 123731 273790 123737 274266
rect 123771 273790 123777 274266
rect 123889 274266 123935 274278
rect 123889 274044 123895 274266
rect 123731 273778 123777 273790
rect 123850 273790 123895 274044
rect 123929 273790 123935 274266
rect 123850 273778 123935 273790
rect 124147 274266 124193 274278
rect 124147 273790 124153 274266
rect 124187 273790 124193 274266
rect 124147 273778 124193 273790
rect 124305 274266 124351 274278
rect 124305 273790 124311 274266
rect 124345 273790 124351 274266
rect 124305 273778 124351 273790
rect 124563 274266 124609 274278
rect 124563 273790 124569 274266
rect 124603 273790 124609 274266
rect 124563 273778 124609 273790
rect 122281 273740 122473 273746
rect 122281 273706 122293 273740
rect 122461 273706 122473 273740
rect 122281 273700 122473 273706
rect 121803 273543 121934 273605
rect 121535 273481 121581 273493
rect 122602 273468 122652 273778
rect 122697 273740 122889 273746
rect 122697 273706 122709 273740
rect 122877 273706 122889 273740
rect 122697 273700 122889 273706
rect 123018 273477 123068 273778
rect 123113 273740 123305 273746
rect 123113 273706 123125 273740
rect 123293 273706 123305 273740
rect 123113 273700 123305 273706
rect 123434 273477 123484 273778
rect 123529 273740 123721 273746
rect 123529 273706 123541 273740
rect 123709 273706 123721 273740
rect 123529 273700 123721 273706
rect 122602 273451 122755 273468
rect 117461 273420 117549 273432
rect 115862 273390 116362 273420
rect 115862 273384 117205 273390
rect 115862 273379 116117 273384
rect 116105 273350 116117 273379
rect 117193 273350 117205 273384
rect 116105 273344 117205 273350
rect 115589 273297 115635 273309
rect 115809 273312 115881 273328
rect 114657 273281 114857 273287
rect 114657 273247 114669 273281
rect 114845 273247 114857 273281
rect 114657 273241 114857 273247
rect 115348 273281 115548 273287
rect 115348 273247 115360 273281
rect 115536 273247 115548 273281
rect 115348 273241 115548 273247
rect 114324 273197 114396 273229
rect 115809 273229 115828 273312
rect 115863 273229 115881 273312
rect 114843 273197 115030 273212
rect 114324 273152 114781 273197
rect 112874 273036 112922 273126
rect 113000 273086 114100 273092
rect 113000 273052 113012 273086
rect 114088 273052 114100 273086
rect 113000 273046 114100 273052
rect 114178 273036 114226 273126
rect 114737 273097 114781 273152
rect 114843 273145 114868 273197
rect 114966 273145 115030 273197
rect 114843 273127 115030 273145
rect 115175 273197 115362 273212
rect 115809 273197 115881 273229
rect 115175 273145 115239 273197
rect 115337 273145 115362 273197
rect 115175 273127 115362 273145
rect 115424 273152 115881 273197
rect 115979 273322 116073 273334
rect 115979 273274 116033 273322
rect 116067 273274 116073 273322
rect 115979 273262 116073 273274
rect 117237 273322 117331 273334
rect 117237 273274 117243 273322
rect 117277 273274 117331 273322
rect 117237 273262 117331 273274
rect 115979 273170 116027 273262
rect 116105 273246 117205 273252
rect 116105 273212 116117 273246
rect 117193 273212 117205 273246
rect 116105 273206 117205 273212
rect 117283 273170 117331 273262
rect 115424 273097 115468 273152
rect 115979 273126 117331 273170
rect 114657 273091 114857 273097
rect 114657 273057 114669 273091
rect 114845 273057 114857 273091
rect 114657 273051 114857 273057
rect 115348 273091 115548 273097
rect 115348 273057 115360 273091
rect 115536 273057 115548 273091
rect 115348 273051 115548 273057
rect 112874 273024 112968 273036
rect 112874 272976 112928 273024
rect 112962 272976 112968 273024
rect 112874 272964 112968 272976
rect 114132 273024 114226 273036
rect 114132 272976 114138 273024
rect 114172 272976 114226 273024
rect 114132 272964 114226 272976
rect 114570 273029 114616 273041
rect 111524 272904 112624 272910
rect 111524 272870 111536 272904
rect 112612 272870 112624 272904
rect 111524 272866 112624 272870
rect 112874 272870 112922 272964
rect 114327 272959 114395 272960
rect 114570 272959 114576 273029
rect 113000 272948 114100 272954
rect 113000 272914 113012 272948
rect 114088 272914 114100 272948
rect 113000 272908 114100 272914
rect 114327 272901 114576 272959
rect 114610 272901 114616 273029
rect 114327 272899 114616 272901
rect 114327 272870 114395 272899
rect 114570 272889 114616 272899
rect 114898 273029 114944 273041
rect 114898 272901 114904 273029
rect 114938 272901 114944 273029
rect 114898 272889 114944 272901
rect 115261 273029 115307 273041
rect 115261 272901 115267 273029
rect 115301 272901 115307 273029
rect 115261 272889 115307 272901
rect 115589 273029 115635 273041
rect 115589 272901 115595 273029
rect 115629 272959 115635 273029
rect 115979 273036 116027 273126
rect 116105 273086 117205 273092
rect 116105 273052 116117 273086
rect 117193 273052 117205 273086
rect 116105 273046 117205 273052
rect 117283 273036 117331 273126
rect 115979 273024 116073 273036
rect 115979 272976 116033 273024
rect 116067 272976 116073 273024
rect 115979 272964 116073 272976
rect 117237 273024 117331 273036
rect 117237 272976 117243 273024
rect 117277 272976 117331 273024
rect 117237 272964 117331 272976
rect 115810 272959 115878 272960
rect 115629 272901 115878 272959
rect 116105 272948 117205 272954
rect 116105 272914 116117 272948
rect 117193 272914 117205 272948
rect 116105 272908 117205 272914
rect 115589 272899 115878 272901
rect 115589 272889 115635 272899
rect 112874 272866 114395 272870
rect 111524 272864 114395 272866
rect 112044 272830 114395 272864
rect 114657 272873 114857 272879
rect 114657 272839 114669 272873
rect 114845 272839 114857 272873
rect 114657 272833 114857 272839
rect 115348 272873 115548 272879
rect 115348 272839 115360 272873
rect 115536 272839 115548 272873
rect 115348 272833 115548 272839
rect 115810 272870 115878 272899
rect 117283 272870 117331 272964
rect 117461 273292 117509 273420
rect 117543 273292 117549 273420
rect 117461 273280 117549 273292
rect 118713 273420 118801 273432
rect 118713 273292 118719 273420
rect 118753 273292 118801 273420
rect 118713 273280 118801 273292
rect 117461 273072 117503 273280
rect 117581 273264 118681 273270
rect 117581 273230 117593 273264
rect 118669 273230 118681 273264
rect 117581 273224 118681 273230
rect 117581 273122 118681 273128
rect 117581 273088 117593 273122
rect 118669 273088 118681 273122
rect 117581 273082 118681 273088
rect 118759 273072 118801 273280
rect 120433 273434 120825 273440
rect 120433 273400 120445 273434
rect 120813 273400 120825 273434
rect 120433 273278 120825 273400
rect 120433 273244 120445 273278
rect 120813 273244 120825 273278
rect 120433 273238 120825 273244
rect 121133 273434 121525 273440
rect 121133 273400 121145 273434
rect 121513 273400 121525 273434
rect 121133 273278 121525 273400
rect 122602 273395 122640 273451
rect 122717 273395 122755 273451
rect 122602 273371 122755 273395
rect 123018 273420 123484 273477
rect 123850 273468 123900 273778
rect 123945 273740 124137 273746
rect 123945 273706 123957 273740
rect 124125 273706 124137 273740
rect 123945 273700 124137 273706
rect 124361 273740 124553 273746
rect 124361 273706 124373 273740
rect 124541 273706 124553 273740
rect 124361 273700 124553 273706
rect 124865 273477 124921 274397
rect 123747 273451 123900 273468
rect 123018 273320 123689 273420
rect 123747 273395 123785 273451
rect 123862 273395 123900 273451
rect 123747 273371 123900 273395
rect 124396 273399 124921 273477
rect 121133 273244 121145 273278
rect 121513 273244 121525 273278
rect 121133 273238 121525 273244
rect 117461 273060 117549 273072
rect 117461 272932 117509 273060
rect 117543 272932 117549 273060
rect 117461 272920 117549 272932
rect 118713 273060 118801 273072
rect 118713 272932 118719 273060
rect 118753 272932 118801 273060
rect 118713 272920 118801 272932
rect 120377 273185 120423 273197
rect 115810 272866 117331 272870
rect 117581 272904 118681 272910
rect 117581 272870 117593 272904
rect 118669 272870 118681 272904
rect 117581 272866 118681 272870
rect 115810 272864 118681 272866
rect 112719 272788 112924 272830
rect 113982 272756 114266 272766
rect 114724 272756 114783 272833
rect 113982 272753 114783 272756
rect 113982 272684 114010 272753
rect 114237 272684 114783 272753
rect 113982 272667 114783 272684
rect 114928 272793 115275 272825
rect 113982 272666 114266 272667
rect 114928 272540 114982 272793
rect 109394 272507 109556 272513
rect 109394 272473 109456 272507
rect 109494 272473 109556 272507
rect 109394 272467 109556 272473
rect 109388 272414 109434 272426
rect 106985 272157 108373 272215
rect 106985 272043 107187 272157
rect 107463 272151 108075 272157
rect 107463 272117 107475 272151
rect 108063 272117 108075 272151
rect 107463 272111 108075 272117
rect 106985 272009 106997 272043
rect 107175 272009 107187 272043
rect 106985 272003 107187 272009
rect 107407 272067 107453 272079
rect 107407 271971 107413 272067
rect 106929 271959 106975 271971
rect 106929 271819 106935 271959
rect 106969 271819 106975 271959
rect 106929 271807 106975 271819
rect 107197 271959 107413 271971
rect 107197 271819 107203 271959
rect 107237 271953 107413 271959
rect 107237 271829 107275 271953
rect 107377 271829 107413 271953
rect 107237 271819 107413 271829
rect 107197 271807 107413 271819
rect 106951 271769 107187 271775
rect 106951 271735 106997 271769
rect 107175 271735 107187 271769
rect 107407 271747 107413 271807
rect 107447 271747 107453 272067
rect 107407 271735 107453 271747
rect 108085 272067 108131 272079
rect 108085 271747 108091 272067
rect 108125 271985 108131 272067
rect 108243 271985 108373 272157
rect 108595 272088 108841 272113
rect 109388 272088 109394 272414
rect 108595 272083 109394 272088
rect 108595 272021 108641 272083
rect 108841 272021 109394 272083
rect 108595 272010 109394 272021
rect 108595 271995 108841 272010
rect 108125 271821 108373 271985
rect 108125 271747 108131 271821
rect 108085 271735 108131 271747
rect 106951 271637 107187 271735
rect 107463 271697 108075 271703
rect 107463 271663 107475 271697
rect 108063 271663 108075 271697
rect 107463 271637 108075 271663
rect 106951 271587 108075 271637
rect 106951 271485 107027 271587
rect 107463 271541 108075 271587
rect 108265 271659 108373 271821
rect 108265 271611 108507 271659
rect 108265 271541 108373 271611
rect 107173 271535 108373 271541
rect 107173 271501 107185 271535
rect 108361 271501 108373 271535
rect 107173 271495 108373 271501
rect 108465 271485 108507 271611
rect 106951 271473 107141 271485
rect 106951 271327 107049 271473
rect 107135 271327 107141 271473
rect 106951 271315 107141 271327
rect 108405 271473 108507 271485
rect 108405 271327 108411 271473
rect 108497 271327 108507 271473
rect 108405 271315 108507 271327
rect 106951 271313 107039 271315
rect 106951 271115 106965 271313
rect 107021 271213 107039 271313
rect 107173 271299 108373 271305
rect 107173 271265 107185 271299
rect 108361 271265 108373 271299
rect 107173 271259 108373 271265
rect 108103 271217 108697 271259
rect 107021 271177 107229 271213
rect 107021 271115 107039 271177
rect 107173 271171 107229 271177
rect 107173 271165 108373 271171
rect 107173 271131 107185 271165
rect 108361 271131 108373 271165
rect 107173 271125 108373 271131
rect 106951 271103 107141 271115
rect 106951 270957 107049 271103
rect 107135 270957 107141 271103
rect 106951 270945 107141 270957
rect 108405 271103 108507 271115
rect 108405 270957 108411 271103
rect 108497 270957 108507 271103
rect 108405 270945 108507 270957
rect 108551 271029 108697 271217
rect 108551 271005 109106 271029
rect 107173 270929 108373 270935
rect 107173 270895 107185 270929
rect 108361 270895 108373 270929
rect 107173 270891 108373 270895
rect 108551 270891 108976 271005
rect 107173 270889 108976 270891
rect 108103 270837 108976 270889
rect 109077 270837 109106 271005
rect 108103 270811 109106 270837
rect 108776 270099 109055 270811
rect 109388 270718 109394 272010
rect 109428 270718 109434 272414
rect 109388 270706 109434 270718
rect 109516 272414 109562 272426
rect 109516 270718 109522 272414
rect 109556 270718 109562 272414
rect 109516 270706 109562 270718
rect 110973 272417 114982 272540
rect 115228 272417 115275 272793
rect 115422 272756 115481 272833
rect 115810 272830 118161 272864
rect 117281 272788 117486 272830
rect 115939 272756 116223 272766
rect 115422 272753 116223 272756
rect 115422 272684 115968 272753
rect 116195 272684 116223 272753
rect 120377 272709 120383 273185
rect 120417 272709 120423 273185
rect 120377 272697 120423 272709
rect 120835 273185 120881 273197
rect 120835 272709 120841 273185
rect 120875 273008 120881 273185
rect 121077 273185 121123 273197
rect 121077 273008 121083 273185
rect 120875 273000 121083 273008
rect 120875 272881 120958 273000
rect 120875 272709 120881 272881
rect 120835 272697 120881 272709
rect 120953 272718 120958 272881
rect 121013 272881 121083 273000
rect 121013 272718 121018 272881
rect 115422 272667 116223 272684
rect 115939 272666 116223 272667
rect 120433 272650 120825 272656
rect 120433 272616 120445 272650
rect 120813 272616 120825 272650
rect 120433 272494 120825 272616
rect 120433 272460 120445 272494
rect 120813 272460 120825 272494
rect 120433 272454 120825 272460
rect 110973 272309 115275 272417
rect 120377 272401 120423 272413
rect 110973 272303 115138 272309
rect 109444 270659 109506 270665
rect 109394 270625 109456 270659
rect 109494 270625 109556 270659
rect 109394 270609 109556 270625
rect 105964 269820 109055 270099
rect 110973 266766 111559 272303
rect 113799 272014 114103 272303
rect 116590 272226 118192 272248
rect 116590 272129 116628 272226
rect 115787 272127 116628 272129
rect 118134 272129 118192 272226
rect 118134 272127 118629 272129
rect 115787 272096 118629 272127
rect 113799 272003 113840 272014
rect 113800 271699 113840 272003
rect 114065 272003 114103 272014
rect 114761 272016 115601 272048
rect 114761 272012 115017 272016
rect 114065 271699 114102 272003
rect 114761 271817 114825 272012
rect 115559 271918 115601 272016
rect 115527 271817 115601 271918
rect 114761 271763 115601 271817
rect 115787 271924 115829 272096
rect 115885 271996 116037 272002
rect 115885 271962 115897 271996
rect 116025 271962 116037 271996
rect 115885 271956 116037 271962
rect 116187 271924 116229 272096
rect 116285 271996 116437 272002
rect 116285 271962 116297 271996
rect 116425 271962 116437 271996
rect 116285 271956 116437 271962
rect 116587 271924 116629 272096
rect 116685 271996 116837 272002
rect 116685 271962 116697 271996
rect 116825 271962 116837 271996
rect 116685 271956 116837 271962
rect 116987 271924 117029 272096
rect 117085 271996 117237 272002
rect 117085 271962 117097 271996
rect 117225 271962 117237 271996
rect 117085 271956 117237 271962
rect 117387 271924 117429 272096
rect 117485 271996 117637 272002
rect 117485 271962 117497 271996
rect 117625 271962 117637 271996
rect 117485 271956 117637 271962
rect 117787 271924 117829 272096
rect 117885 271996 118037 272002
rect 117885 271962 117897 271996
rect 118025 271962 118037 271996
rect 117885 271956 118037 271962
rect 118187 271924 118229 272096
rect 118285 271996 118437 272002
rect 118285 271962 118297 271996
rect 118425 271962 118437 271996
rect 118285 271956 118437 271962
rect 118587 271924 118629 272096
rect 118685 271996 118837 272002
rect 118685 271962 118697 271996
rect 118825 271962 118837 271996
rect 118685 271956 118837 271962
rect 120377 271925 120383 272401
rect 120417 271925 120423 272401
rect 115787 271912 115875 271924
rect 113800 271668 114102 271699
rect 113068 271629 113461 271643
rect 113068 271540 113091 271629
rect 113431 271540 113461 271629
rect 112790 271501 113726 271540
rect 112582 271387 112734 271393
rect 112582 271353 112594 271387
rect 112722 271353 112734 271387
rect 112582 271347 112734 271353
rect 112790 271306 112840 271501
rect 112982 271387 113134 271393
rect 112982 271353 112994 271387
rect 113122 271353 113134 271387
rect 112982 271347 113134 271353
rect 113233 271306 113283 271501
rect 113382 271387 113534 271393
rect 113382 271353 113394 271387
rect 113522 271353 113534 271387
rect 113382 271347 113534 271353
rect 113676 271306 113726 271501
rect 113782 271387 114490 271393
rect 113782 271353 113794 271387
rect 113922 271353 114490 271387
rect 115091 271364 115154 271763
rect 113782 271347 114490 271353
rect 113900 271346 114490 271347
rect 112484 271294 112572 271306
rect 112484 271118 112532 271294
rect 112566 271118 112572 271294
rect 112484 271106 112572 271118
rect 112744 271294 112840 271306
rect 112744 271118 112750 271294
rect 112784 271118 112840 271294
rect 112744 271106 112840 271118
rect 112884 271294 112972 271306
rect 112884 271118 112932 271294
rect 112966 271118 112972 271294
rect 112884 271106 112972 271118
rect 113144 271294 113372 271306
rect 113144 271118 113150 271294
rect 113184 271247 113332 271294
rect 113184 271118 113190 271247
rect 113144 271106 113190 271118
rect 113326 271118 113332 271247
rect 113366 271118 113372 271294
rect 113326 271106 113372 271118
rect 113544 271294 113632 271306
rect 113544 271118 113550 271294
rect 113584 271118 113632 271294
rect 113544 271106 113632 271118
rect 113676 271294 113772 271306
rect 113676 271118 113732 271294
rect 113766 271118 113772 271294
rect 113676 271106 113772 271118
rect 113944 271294 114032 271306
rect 113944 271118 113950 271294
rect 113984 271118 114032 271294
rect 114425 271277 114490 271346
rect 114641 271358 115193 271364
rect 114641 271324 114653 271358
rect 114781 271324 115053 271358
rect 115181 271324 115193 271358
rect 114641 271318 115193 271324
rect 114425 271265 114631 271277
rect 114425 271230 114591 271265
rect 113944 271106 114032 271118
rect 112484 270939 112526 271106
rect 112582 271059 112734 271065
rect 112582 271025 112594 271059
rect 112722 271025 112734 271059
rect 112582 271019 112734 271025
rect 112884 270939 112926 271106
rect 112982 271059 113134 271065
rect 112982 271025 112994 271059
rect 113122 271025 113134 271059
rect 112982 271019 113134 271025
rect 113382 271059 113534 271065
rect 113382 271025 113394 271059
rect 113522 271025 113534 271059
rect 113382 271019 113534 271025
rect 113590 270939 113632 271106
rect 113782 271059 113934 271065
rect 113782 271025 113794 271059
rect 113922 271025 113934 271059
rect 113782 271019 113934 271025
rect 113990 270939 114032 271106
rect 112484 270901 114032 270939
rect 114537 271089 114591 271230
rect 114625 271089 114631 271265
rect 114537 271077 114631 271089
rect 114803 271265 114849 271277
rect 114803 271089 114809 271265
rect 114843 271089 114849 271265
rect 114803 271077 114849 271089
rect 114985 271265 115031 271277
rect 114985 271089 114991 271265
rect 115025 271089 115031 271265
rect 114985 271077 115031 271089
rect 115203 271265 115297 271277
rect 115203 271089 115209 271265
rect 115243 271089 115297 271265
rect 115203 271077 115297 271089
rect 114537 270909 114585 271077
rect 114641 271030 114793 271036
rect 114641 270996 114653 271030
rect 114781 270996 114793 271030
rect 114641 270990 114793 270996
rect 115041 271030 115193 271036
rect 115041 270996 115053 271030
rect 115181 270996 115193 271030
rect 115041 270990 115193 270996
rect 115249 270909 115297 271077
rect 112676 270715 112792 270901
rect 114537 270869 115297 270909
rect 112194 270671 113508 270715
rect 112194 270446 112267 270671
rect 113449 270446 113508 270671
rect 114050 270673 114542 270693
rect 114050 270576 114086 270673
rect 114501 270657 114542 270673
rect 114850 270657 114976 270869
rect 115787 270836 115835 271912
rect 115869 270836 115875 271912
rect 115787 270824 115875 270836
rect 116047 271912 116135 271924
rect 116047 270836 116053 271912
rect 116087 270836 116135 271912
rect 116047 270824 116135 270836
rect 116187 271912 116275 271924
rect 116187 270836 116235 271912
rect 116269 270836 116275 271912
rect 116187 270824 116275 270836
rect 116447 271912 116535 271924
rect 116447 270836 116453 271912
rect 116487 270836 116535 271912
rect 116447 270824 116535 270836
rect 116587 271912 116675 271924
rect 116587 270836 116635 271912
rect 116669 270836 116675 271912
rect 116587 270824 116675 270836
rect 116847 271912 116935 271924
rect 116847 270836 116853 271912
rect 116887 270836 116935 271912
rect 116847 270824 116935 270836
rect 116987 271912 117075 271924
rect 116987 270836 117035 271912
rect 117069 270836 117075 271912
rect 116987 270824 117075 270836
rect 117247 271912 117335 271924
rect 117247 270836 117253 271912
rect 117287 270836 117335 271912
rect 117247 270824 117335 270836
rect 117387 271912 117475 271924
rect 117387 270836 117435 271912
rect 117469 270836 117475 271912
rect 117387 270824 117475 270836
rect 117647 271912 117735 271924
rect 117647 270836 117653 271912
rect 117687 270836 117735 271912
rect 117647 270824 117735 270836
rect 117787 271912 117875 271924
rect 117787 270836 117835 271912
rect 117869 270836 117875 271912
rect 117787 270824 117875 270836
rect 118047 271912 118135 271924
rect 118047 270836 118053 271912
rect 118087 270836 118135 271912
rect 118047 270824 118135 270836
rect 118187 271912 118275 271924
rect 118187 270836 118235 271912
rect 118269 270836 118275 271912
rect 118187 270824 118275 270836
rect 118447 271912 118535 271924
rect 118447 270836 118453 271912
rect 118487 270836 118535 271912
rect 118447 270824 118535 270836
rect 118587 271912 118675 271924
rect 118587 270836 118635 271912
rect 118669 270836 118675 271912
rect 118587 270824 118675 270836
rect 118847 271912 118935 271924
rect 120377 271913 120423 271925
rect 120835 272401 120881 272413
rect 120835 271925 120841 272401
rect 120875 272224 120881 272401
rect 120953 272224 121018 272718
rect 121077 272709 121083 272881
rect 121117 272709 121123 273185
rect 121077 272697 121123 272709
rect 121535 273185 121624 273197
rect 121535 272709 121541 273185
rect 121575 272709 121624 273185
rect 121535 272697 121624 272709
rect 121133 272650 121525 272656
rect 121133 272616 121145 272650
rect 121513 272616 121525 272650
rect 121133 272494 121525 272616
rect 121133 272460 121145 272494
rect 121513 272460 121525 272494
rect 121133 272454 121525 272460
rect 121581 272413 121624 272697
rect 121796 273059 123438 273127
rect 121077 272401 121123 272413
rect 121077 272224 121083 272401
rect 120875 272097 121083 272224
rect 120875 271925 120881 272097
rect 120835 271913 120881 271925
rect 118847 270836 118853 271912
rect 118887 270836 118935 271912
rect 120433 271866 120825 271872
rect 120433 271832 120445 271866
rect 120813 271832 120825 271866
rect 120433 271710 120825 271832
rect 120433 271676 120445 271710
rect 120813 271676 120825 271710
rect 120433 271670 120825 271676
rect 120377 271617 120423 271629
rect 120377 271141 120383 271617
rect 120417 271141 120423 271617
rect 120377 271129 120423 271141
rect 120835 271617 120881 271629
rect 120835 271141 120841 271617
rect 120875 271440 120881 271617
rect 120953 271440 121018 272097
rect 121077 271925 121083 272097
rect 121117 271925 121123 272401
rect 121077 271913 121123 271925
rect 121535 272401 121677 272413
rect 121535 271925 121541 272401
rect 121575 272340 121677 272401
rect 121575 271925 121605 272340
rect 121535 271913 121605 271925
rect 121133 271866 121525 271872
rect 121133 271832 121145 271866
rect 121513 271832 121525 271866
rect 121133 271710 121525 271832
rect 121133 271676 121145 271710
rect 121513 271676 121525 271710
rect 121133 271670 121525 271676
rect 121581 271629 121605 271913
rect 121077 271617 121123 271629
rect 121077 271440 121083 271617
rect 120875 271313 121083 271440
rect 120875 271141 120881 271313
rect 120835 271129 120881 271141
rect 120433 271082 120825 271088
rect 120433 271048 120445 271082
rect 120813 271048 120825 271082
rect 120433 270926 120825 271048
rect 120433 270892 120445 270926
rect 120813 270892 120825 270926
rect 120433 270886 120825 270892
rect 118847 270824 118935 270836
rect 115885 270786 116037 270792
rect 115885 270752 115897 270786
rect 116025 270752 116037 270786
rect 115885 270746 116037 270752
rect 114501 270617 114976 270657
rect 116093 270621 116135 270824
rect 116285 270786 116437 270792
rect 116285 270752 116297 270786
rect 116425 270752 116437 270786
rect 116285 270746 116437 270752
rect 116493 270621 116535 270824
rect 116685 270786 116837 270792
rect 116685 270752 116697 270786
rect 116825 270752 116837 270786
rect 116685 270746 116837 270752
rect 116893 270621 116935 270824
rect 117085 270786 117237 270792
rect 117085 270752 117097 270786
rect 117225 270752 117237 270786
rect 117085 270746 117237 270752
rect 117293 270621 117335 270824
rect 117485 270786 117637 270792
rect 117485 270752 117497 270786
rect 117625 270752 117637 270786
rect 117485 270746 117637 270752
rect 117693 270621 117735 270824
rect 117885 270786 118037 270792
rect 117885 270752 117897 270786
rect 118025 270752 118037 270786
rect 117885 270746 118037 270752
rect 118093 270621 118135 270824
rect 118285 270786 118437 270792
rect 118285 270752 118297 270786
rect 118425 270752 118437 270786
rect 118285 270746 118437 270752
rect 118493 270621 118535 270824
rect 118685 270786 118837 270792
rect 118685 270752 118697 270786
rect 118825 270752 118837 270786
rect 118685 270746 118837 270752
rect 118893 270621 118935 270824
rect 116093 270617 118935 270621
rect 114501 270588 118935 270617
rect 120377 270833 120423 270845
rect 114501 270587 116771 270588
rect 114501 270586 114877 270587
rect 114501 270576 114542 270586
rect 114050 270545 114542 270576
rect 112194 270429 113508 270446
rect 112194 270399 118508 270429
rect 112466 270396 118508 270399
rect 112466 270224 112508 270396
rect 112564 270296 112716 270302
rect 112564 270262 112576 270296
rect 112704 270262 112716 270296
rect 112564 270256 112716 270262
rect 112866 270224 112908 270396
rect 112964 270296 113116 270302
rect 112964 270262 112976 270296
rect 113104 270262 113116 270296
rect 112964 270256 113116 270262
rect 113266 270224 113308 270396
rect 113364 270296 113516 270302
rect 113364 270262 113376 270296
rect 113504 270262 113516 270296
rect 113364 270256 113516 270262
rect 113666 270224 113708 270396
rect 113764 270296 113916 270302
rect 113764 270262 113776 270296
rect 113904 270262 113916 270296
rect 113764 270256 113916 270262
rect 114066 270224 114108 270396
rect 114164 270296 114316 270302
rect 114164 270262 114176 270296
rect 114304 270262 114316 270296
rect 114164 270256 114316 270262
rect 114466 270224 114508 270396
rect 114564 270296 114716 270302
rect 114564 270262 114576 270296
rect 114704 270262 114716 270296
rect 114564 270256 114716 270262
rect 114866 270224 114908 270396
rect 114964 270296 115116 270302
rect 114964 270262 114976 270296
rect 115104 270262 115116 270296
rect 114964 270256 115116 270262
rect 115266 270224 115308 270396
rect 115364 270296 115516 270302
rect 115364 270262 115376 270296
rect 115504 270262 115516 270296
rect 115364 270256 115516 270262
rect 115666 270224 115708 270396
rect 115764 270296 115916 270302
rect 115764 270262 115776 270296
rect 115904 270262 115916 270296
rect 115764 270256 115916 270262
rect 116066 270224 116108 270396
rect 116164 270296 116316 270302
rect 116164 270262 116176 270296
rect 116304 270262 116316 270296
rect 116164 270256 116316 270262
rect 116466 270224 116508 270396
rect 116564 270296 116716 270302
rect 116564 270262 116576 270296
rect 116704 270262 116716 270296
rect 116564 270256 116716 270262
rect 116866 270224 116908 270396
rect 116964 270296 117116 270302
rect 116964 270262 116976 270296
rect 117104 270262 117116 270296
rect 116964 270256 117116 270262
rect 117266 270224 117308 270396
rect 117364 270296 117516 270302
rect 117364 270262 117376 270296
rect 117504 270262 117516 270296
rect 117364 270256 117516 270262
rect 117666 270224 117708 270396
rect 117764 270296 117916 270302
rect 117764 270262 117776 270296
rect 117904 270262 117916 270296
rect 117764 270256 117916 270262
rect 118066 270224 118108 270396
rect 118164 270296 118316 270302
rect 118164 270262 118176 270296
rect 118304 270262 118316 270296
rect 118164 270256 118316 270262
rect 118466 270224 118508 270396
rect 120377 270357 120383 270833
rect 120417 270357 120423 270833
rect 120377 270345 120423 270357
rect 120835 270833 120881 270845
rect 120835 270357 120841 270833
rect 120875 270656 120881 270833
rect 120953 270656 121018 271313
rect 121077 271141 121083 271313
rect 121117 271141 121123 271617
rect 121077 271129 121123 271141
rect 121535 271617 121605 271629
rect 121535 271141 121541 271617
rect 121575 271141 121605 271617
rect 121535 271129 121605 271141
rect 121133 271082 121525 271088
rect 121133 271048 121145 271082
rect 121513 271048 121525 271082
rect 121133 270926 121525 271048
rect 121133 270892 121145 270926
rect 121513 270892 121525 270926
rect 121133 270886 121525 270892
rect 121581 270845 121605 271129
rect 121077 270833 121123 270845
rect 121077 270656 121083 270833
rect 120875 270529 121083 270656
rect 120875 270357 120881 270529
rect 120835 270345 120881 270357
rect 118564 270296 118716 270302
rect 118564 270262 118576 270296
rect 118704 270262 118716 270296
rect 118564 270256 118716 270262
rect 120433 270298 120825 270304
rect 120433 270264 120445 270298
rect 120813 270264 120825 270298
rect 112466 270212 112554 270224
rect 112466 269136 112514 270212
rect 112548 269136 112554 270212
rect 112466 269124 112554 269136
rect 112726 270212 112814 270224
rect 112726 269136 112732 270212
rect 112766 269136 112814 270212
rect 112726 269124 112814 269136
rect 112866 270212 112954 270224
rect 112866 269136 112914 270212
rect 112948 269136 112954 270212
rect 112866 269124 112954 269136
rect 113126 270212 113214 270224
rect 113126 269136 113132 270212
rect 113166 269136 113214 270212
rect 113126 269124 113214 269136
rect 113266 270212 113354 270224
rect 113266 269136 113314 270212
rect 113348 269136 113354 270212
rect 113266 269124 113354 269136
rect 113526 270212 113614 270224
rect 113526 269136 113532 270212
rect 113566 269136 113614 270212
rect 113526 269124 113614 269136
rect 113666 270212 113754 270224
rect 113666 269136 113714 270212
rect 113748 269136 113754 270212
rect 113666 269124 113754 269136
rect 113926 270212 114014 270224
rect 113926 269136 113932 270212
rect 113966 269136 114014 270212
rect 113926 269124 114014 269136
rect 114066 270212 114154 270224
rect 114066 269136 114114 270212
rect 114148 269136 114154 270212
rect 114066 269124 114154 269136
rect 114326 270212 114414 270224
rect 114326 269136 114332 270212
rect 114366 269136 114414 270212
rect 114326 269124 114414 269136
rect 114466 270212 114554 270224
rect 114466 269136 114514 270212
rect 114548 269136 114554 270212
rect 114466 269124 114554 269136
rect 114726 270212 114814 270224
rect 114726 269136 114732 270212
rect 114766 269136 114814 270212
rect 114726 269124 114814 269136
rect 114866 270212 114954 270224
rect 114866 269136 114914 270212
rect 114948 269136 114954 270212
rect 114866 269124 114954 269136
rect 115126 270212 115214 270224
rect 115126 269136 115132 270212
rect 115166 269136 115214 270212
rect 115126 269124 115214 269136
rect 115266 270212 115354 270224
rect 115266 269136 115314 270212
rect 115348 269136 115354 270212
rect 115266 269124 115354 269136
rect 115526 270212 115614 270224
rect 115526 269136 115532 270212
rect 115566 269136 115614 270212
rect 115526 269124 115614 269136
rect 115666 270212 115754 270224
rect 115666 269136 115714 270212
rect 115748 269136 115754 270212
rect 115666 269124 115754 269136
rect 115926 270212 116014 270224
rect 115926 269136 115932 270212
rect 115966 269136 116014 270212
rect 115926 269124 116014 269136
rect 116066 270212 116154 270224
rect 116066 269136 116114 270212
rect 116148 269136 116154 270212
rect 116066 269124 116154 269136
rect 116326 270212 116414 270224
rect 116326 269136 116332 270212
rect 116366 269136 116414 270212
rect 116326 269124 116414 269136
rect 116466 270212 116554 270224
rect 116466 269136 116514 270212
rect 116548 269136 116554 270212
rect 116466 269124 116554 269136
rect 116726 270212 116814 270224
rect 116726 269136 116732 270212
rect 116766 269136 116814 270212
rect 116726 269124 116814 269136
rect 116866 270212 116954 270224
rect 116866 269136 116914 270212
rect 116948 269136 116954 270212
rect 116866 269124 116954 269136
rect 117126 270212 117214 270224
rect 117126 269136 117132 270212
rect 117166 269136 117214 270212
rect 117126 269124 117214 269136
rect 117266 270212 117354 270224
rect 117266 269136 117314 270212
rect 117348 269136 117354 270212
rect 117266 269124 117354 269136
rect 117526 270212 117614 270224
rect 117526 269136 117532 270212
rect 117566 269136 117614 270212
rect 117526 269124 117614 269136
rect 117666 270212 117754 270224
rect 117666 269136 117714 270212
rect 117748 269136 117754 270212
rect 117666 269124 117754 269136
rect 117926 270212 118014 270224
rect 117926 269136 117932 270212
rect 117966 269136 118014 270212
rect 117926 269124 118014 269136
rect 118066 270212 118154 270224
rect 118066 269136 118114 270212
rect 118148 269136 118154 270212
rect 118066 269124 118154 269136
rect 118326 270212 118414 270224
rect 118326 269136 118332 270212
rect 118366 269136 118414 270212
rect 118326 269124 118414 269136
rect 118466 270212 118554 270224
rect 118466 269136 118514 270212
rect 118548 269136 118554 270212
rect 118466 269124 118554 269136
rect 118726 270212 118814 270224
rect 118726 269136 118732 270212
rect 118766 269136 118814 270212
rect 120433 270142 120825 270264
rect 120433 270108 120445 270142
rect 120813 270108 120825 270142
rect 120433 270102 120825 270108
rect 120377 270049 120423 270061
rect 120377 269573 120383 270049
rect 120417 269573 120423 270049
rect 120377 269561 120423 269573
rect 120835 270049 120881 270061
rect 120835 269573 120841 270049
rect 120875 269872 120881 270049
rect 120953 269872 121018 270529
rect 121077 270357 121083 270529
rect 121117 270357 121123 270833
rect 121077 270345 121123 270357
rect 121535 270833 121605 270845
rect 121535 270357 121541 270833
rect 121575 270428 121605 270833
rect 121657 270428 121677 272340
rect 121575 270357 121677 270428
rect 121535 270345 121677 270357
rect 121133 270298 121525 270304
rect 121133 270264 121145 270298
rect 121513 270264 121525 270298
rect 121133 270142 121525 270264
rect 121133 270108 121145 270142
rect 121513 270108 121525 270142
rect 121133 270102 121525 270108
rect 121581 270061 121624 270345
rect 121077 270049 121123 270061
rect 121077 269872 121083 270049
rect 120875 269745 121083 269872
rect 120875 269573 120881 269745
rect 120835 269561 120881 269573
rect 121077 269573 121083 269745
rect 121117 269573 121123 270049
rect 121077 269561 121123 269573
rect 121535 270049 121624 270061
rect 121535 269573 121541 270049
rect 121575 269573 121624 270049
rect 121535 269561 121624 269573
rect 120433 269514 120825 269520
rect 120433 269480 120445 269514
rect 120813 269480 120825 269514
rect 121133 269514 121525 269520
rect 121133 269496 121145 269514
rect 120433 269474 120825 269480
rect 121132 269480 121145 269496
rect 121513 269496 121525 269514
rect 121796 269496 121864 273059
rect 122129 272894 122521 272900
rect 122129 272860 122141 272894
rect 122509 272860 122521 272894
rect 122129 272854 122521 272860
rect 122829 272894 123221 272900
rect 122829 272860 122841 272894
rect 123209 272860 123221 272894
rect 122829 272854 123221 272860
rect 122073 272801 122119 272813
rect 122073 272725 122079 272801
rect 122113 272725 122119 272801
rect 122073 272713 122119 272725
rect 122531 272801 122577 272813
rect 122531 272725 122537 272801
rect 122571 272725 122577 272801
rect 122531 272713 122577 272725
rect 122773 272801 122819 272813
rect 122773 272725 122779 272801
rect 122813 272725 122819 272801
rect 122773 272713 122819 272725
rect 123231 272801 123277 272813
rect 123231 272725 123237 272801
rect 123271 272725 123277 272801
rect 123231 272713 123277 272725
rect 122129 272666 122521 272672
rect 122129 272632 122141 272666
rect 122509 272632 122521 272666
rect 122129 272626 122521 272632
rect 122829 272666 123221 272672
rect 122829 272632 122841 272666
rect 123209 272632 123221 272666
rect 123368 272656 123438 273059
rect 122829 272626 123221 272632
rect 123333 272626 123462 272656
rect 121513 269480 121864 269496
rect 121132 269436 121864 269480
rect 121991 272510 122521 272516
rect 121991 272476 122141 272510
rect 122509 272476 122521 272510
rect 121991 272470 122521 272476
rect 122829 272510 123221 272516
rect 122829 272476 122841 272510
rect 123209 272476 123221 272510
rect 122829 272470 123221 272476
rect 121991 271888 122023 272470
rect 123333 272446 123355 272626
rect 123444 272446 123462 272626
rect 122073 272417 122119 272429
rect 122073 271941 122079 272417
rect 122113 271941 122119 272417
rect 122073 271929 122119 271941
rect 122531 272417 122577 272429
rect 122531 271941 122537 272417
rect 122571 272235 122577 272417
rect 122773 272417 122819 272429
rect 122773 272235 122779 272417
rect 122571 272214 122779 272235
rect 122571 272150 122654 272214
rect 122710 272150 122779 272214
rect 122571 272128 122779 272150
rect 122571 271941 122577 272128
rect 122531 271929 122577 271941
rect 121991 271882 122521 271888
rect 121991 271848 122141 271882
rect 122509 271848 122521 271882
rect 121991 271842 122521 271848
rect 121991 271732 122023 271842
rect 121991 271726 122521 271732
rect 121991 271692 122141 271726
rect 122509 271692 122521 271726
rect 121991 271686 122521 271692
rect 121991 271104 122023 271686
rect 122073 271633 122119 271645
rect 122073 271157 122079 271633
rect 122113 271157 122119 271633
rect 122073 271145 122119 271157
rect 122531 271633 122577 271645
rect 122531 271157 122537 271633
rect 122571 271157 122577 271633
rect 122531 271145 122577 271157
rect 121991 271098 122521 271104
rect 121991 271064 122141 271098
rect 122509 271064 122521 271098
rect 121991 271058 122521 271064
rect 121991 270948 122023 271058
rect 121991 270942 122521 270948
rect 121991 270908 122141 270942
rect 122509 270908 122521 270942
rect 121991 270902 122521 270908
rect 121991 270320 122023 270902
rect 122073 270849 122119 270861
rect 122073 270373 122079 270849
rect 122113 270373 122119 270849
rect 122073 270361 122119 270373
rect 122531 270849 122577 270861
rect 122531 270373 122537 270849
rect 122571 270373 122577 270849
rect 122531 270361 122577 270373
rect 121991 270314 122521 270320
rect 121991 270280 122141 270314
rect 122509 270280 122521 270314
rect 121991 270274 122521 270280
rect 121991 270164 122023 270274
rect 121991 270158 122521 270164
rect 121991 270124 122141 270158
rect 122509 270124 122521 270158
rect 121991 270118 122521 270124
rect 121991 269536 122023 270118
rect 122073 270065 122119 270077
rect 122073 269589 122079 270065
rect 122113 269589 122119 270065
rect 122073 269577 122119 269589
rect 122531 270065 122577 270077
rect 122531 269589 122537 270065
rect 122571 269874 122577 270065
rect 122646 269874 122724 272128
rect 122773 271941 122779 272128
rect 122813 271941 122819 272417
rect 122773 271929 122819 271941
rect 123231 272417 123277 272429
rect 123333 272427 123462 272446
rect 123231 271941 123237 272417
rect 123271 272231 123277 272417
rect 123362 272231 123476 272233
rect 123271 272200 123476 272231
rect 123271 272125 123380 272200
rect 123271 272124 123329 272125
rect 123271 271941 123277 272124
rect 123362 272040 123380 272125
rect 123463 272194 123476 272200
rect 123595 272194 123689 273320
rect 124396 273110 124462 273399
rect 123463 272083 123689 272194
rect 123774 273024 124462 273110
rect 124634 273042 124956 273071
rect 123463 272040 123476 272083
rect 123362 272007 123476 272040
rect 123231 271929 123277 271941
rect 122829 271882 123221 271888
rect 122829 271848 122841 271882
rect 123209 271848 123221 271882
rect 122829 271726 123221 271848
rect 122829 271692 122841 271726
rect 123209 271692 123221 271726
rect 122829 271686 123221 271692
rect 122773 271633 122819 271645
rect 122773 271157 122779 271633
rect 122813 271157 122819 271633
rect 122773 271145 122819 271157
rect 123231 271633 123337 271645
rect 123231 271157 123237 271633
rect 123271 271157 123337 271633
rect 123231 271145 123337 271157
rect 122829 271098 123221 271104
rect 122829 271064 122841 271098
rect 123209 271064 123221 271098
rect 122829 270942 123221 271064
rect 122829 270908 122841 270942
rect 123209 270908 123221 270942
rect 122829 270902 123221 270908
rect 123277 271065 123337 271145
rect 123774 271440 123842 273024
rect 124634 272915 124666 273042
rect 123930 272845 124666 272915
rect 124931 272845 124956 273042
rect 123930 272816 124956 272845
rect 123930 271856 123993 272816
rect 124634 272811 124956 272816
rect 124192 272566 124692 272572
rect 124192 272532 124204 272566
rect 124680 272532 124692 272566
rect 124192 272526 124692 272532
rect 124114 272504 124160 272516
rect 124114 272336 124120 272504
rect 124154 272336 124160 272504
rect 124114 272324 124160 272336
rect 124724 272504 124770 272516
rect 124724 272336 124730 272504
rect 124764 272336 124770 272504
rect 124724 272320 124770 272336
rect 124192 272308 124692 272314
rect 124192 272274 124204 272308
rect 124680 272274 124692 272308
rect 124192 272268 124692 272274
rect 124192 272150 124692 272156
rect 124192 272116 124204 272150
rect 124680 272116 124692 272150
rect 124192 272110 124692 272116
rect 124114 272088 124160 272100
rect 124114 271920 124120 272088
rect 124154 271920 124160 272088
rect 124114 271908 124160 271920
rect 124724 272088 124770 272104
rect 124724 271920 124730 272088
rect 124764 271920 124770 272088
rect 124192 271892 124692 271898
rect 124192 271858 124204 271892
rect 124680 271858 124692 271892
rect 124192 271856 124692 271858
rect 123930 271806 124692 271856
rect 123930 271804 123993 271806
rect 124192 271734 124692 271740
rect 124192 271700 124204 271734
rect 124680 271700 124692 271734
rect 124192 271694 124692 271700
rect 124114 271672 124160 271684
rect 124114 271504 124120 271672
rect 124154 271504 124160 271672
rect 124114 271492 124160 271504
rect 124724 271672 124770 271920
rect 124724 271504 124730 271672
rect 124764 271504 124770 271672
rect 124192 271476 124692 271482
rect 124192 271442 124204 271476
rect 124680 271442 124692 271476
rect 124192 271440 124692 271442
rect 123774 271390 124692 271440
rect 123774 271065 123847 271390
rect 124192 271318 124692 271324
rect 124192 271284 124204 271318
rect 124680 271284 124692 271318
rect 124192 271278 124692 271284
rect 124068 271256 124160 271268
rect 124068 271093 124120 271256
rect 123277 270918 123847 271065
rect 123277 270861 123337 270918
rect 122773 270849 122819 270861
rect 122773 270373 122779 270849
rect 122813 270373 122819 270849
rect 122773 270361 122819 270373
rect 123231 270849 123337 270861
rect 123231 270373 123237 270849
rect 123271 270373 123337 270849
rect 123231 270361 123337 270373
rect 122829 270314 123221 270320
rect 122829 270280 122841 270314
rect 123209 270280 123221 270314
rect 122829 270158 123221 270280
rect 122829 270124 122841 270158
rect 123209 270124 123221 270158
rect 123774 270192 123847 270918
rect 123931 271088 124120 271093
rect 124154 271088 124160 271256
rect 123931 271076 124160 271088
rect 124724 271256 124770 271504
rect 124724 271088 124730 271256
rect 124764 271088 124770 271256
rect 123931 271033 124114 271076
rect 123931 270785 123962 271033
rect 124063 271024 124114 271033
rect 124192 271060 124692 271066
rect 124192 271026 124204 271060
rect 124680 271026 124692 271060
rect 124192 271024 124692 271026
rect 124063 270974 124692 271024
rect 124063 270852 124114 270974
rect 124192 270902 124692 270908
rect 124192 270868 124204 270902
rect 124680 270868 124692 270902
rect 124192 270862 124692 270868
rect 124063 270840 124160 270852
rect 124063 270785 124120 270840
rect 123931 270717 124120 270785
rect 124068 270672 124120 270717
rect 124154 270672 124160 270840
rect 124068 270660 124160 270672
rect 124724 270840 124770 271088
rect 124724 270672 124730 270840
rect 124764 270672 124770 270840
rect 124068 270608 124114 270660
rect 124192 270644 124692 270650
rect 124192 270610 124204 270644
rect 124680 270610 124692 270644
rect 124192 270608 124692 270610
rect 124068 270558 124692 270608
rect 124192 270486 124692 270492
rect 124192 270452 124204 270486
rect 124680 270452 124692 270486
rect 124192 270446 124692 270452
rect 124114 270424 124160 270436
rect 124114 270256 124120 270424
rect 124154 270256 124160 270424
rect 124114 270244 124160 270256
rect 124724 270424 124770 270672
rect 124724 270256 124730 270424
rect 124764 270256 124770 270424
rect 124192 270228 124692 270234
rect 124192 270194 124204 270228
rect 124680 270194 124692 270228
rect 124192 270192 124692 270194
rect 123774 270142 124692 270192
rect 122829 270118 123221 270124
rect 122773 270065 122819 270077
rect 122773 269874 122779 270065
rect 122571 269852 122779 269874
rect 122571 269788 122657 269852
rect 122713 269788 122779 269852
rect 122571 269767 122779 269788
rect 122571 269589 122577 269767
rect 122531 269577 122577 269589
rect 122773 269589 122779 269767
rect 122813 269589 122819 270065
rect 122773 269577 122819 269589
rect 123231 270065 123277 270077
rect 123231 269589 123237 270065
rect 123271 269865 123277 270065
rect 124192 270070 124692 270076
rect 124192 270036 124204 270070
rect 124680 270036 124692 270070
rect 124192 270030 124692 270036
rect 124114 270008 124160 270020
rect 123271 269864 123411 269865
rect 123271 269833 123474 269864
rect 123271 269758 123377 269833
rect 123271 269589 123277 269758
rect 123231 269577 123277 269589
rect 123360 269673 123377 269758
rect 123460 269673 123474 269833
rect 124114 269840 124120 270008
rect 124154 269840 124160 270008
rect 124114 269828 124160 269840
rect 124724 270008 124770 270256
rect 124724 269840 124730 270008
rect 124764 269840 124770 270008
rect 124724 269824 124770 269840
rect 124192 269812 124692 269818
rect 124192 269778 124204 269812
rect 124680 269790 124692 269812
rect 124878 269790 124944 272811
rect 124680 269778 124944 269790
rect 124192 269769 124944 269778
rect 124192 269737 124943 269769
rect 123360 269638 123474 269673
rect 124192 269654 124692 269660
rect 121991 269530 122521 269536
rect 121991 269496 122141 269530
rect 122509 269496 122521 269530
rect 121991 269490 122521 269496
rect 122829 269530 123221 269536
rect 122829 269496 122841 269530
rect 123209 269496 123221 269530
rect 122829 269490 123221 269496
rect 120433 269358 120825 269364
rect 120433 269324 120445 269358
rect 120813 269324 120825 269358
rect 120433 269318 120825 269324
rect 121133 269358 121525 269364
rect 121133 269324 121145 269358
rect 121513 269324 121525 269358
rect 121133 269318 121525 269324
rect 120377 269265 120423 269277
rect 120377 269189 120383 269265
rect 120417 269189 120423 269265
rect 120377 269177 120423 269189
rect 120835 269265 120881 269277
rect 120835 269189 120841 269265
rect 120875 269189 120881 269265
rect 120835 269177 120881 269189
rect 121077 269265 121123 269277
rect 121077 269189 121083 269265
rect 121117 269189 121123 269265
rect 121077 269177 121123 269189
rect 121535 269265 121581 269277
rect 121535 269189 121541 269265
rect 121575 269189 121581 269265
rect 121535 269177 121581 269189
rect 118726 269124 118814 269136
rect 112564 269086 112716 269092
rect 112564 269052 112576 269086
rect 112704 269052 112716 269086
rect 112564 269046 112716 269052
rect 112772 268921 112814 269124
rect 112964 269086 113116 269092
rect 112964 269052 112976 269086
rect 113104 269052 113116 269086
rect 112964 269046 113116 269052
rect 113172 268921 113214 269124
rect 113364 269086 113516 269092
rect 113364 269052 113376 269086
rect 113504 269052 113516 269086
rect 113364 269046 113516 269052
rect 113572 268921 113614 269124
rect 113764 269086 113916 269092
rect 113764 269052 113776 269086
rect 113904 269052 113916 269086
rect 113764 269046 113916 269052
rect 113972 268921 114014 269124
rect 114164 269086 114316 269092
rect 114164 269052 114176 269086
rect 114304 269052 114316 269086
rect 114164 269046 114316 269052
rect 114372 268921 114414 269124
rect 114564 269086 114716 269092
rect 114564 269052 114576 269086
rect 114704 269052 114716 269086
rect 114564 269046 114716 269052
rect 114772 268921 114814 269124
rect 114964 269086 115116 269092
rect 114964 269052 114976 269086
rect 115104 269052 115116 269086
rect 114964 269046 115116 269052
rect 115172 268921 115214 269124
rect 115364 269086 115516 269092
rect 115364 269052 115376 269086
rect 115504 269052 115516 269086
rect 115364 269046 115516 269052
rect 115572 268921 115614 269124
rect 115764 269086 115916 269092
rect 115764 269052 115776 269086
rect 115904 269052 115916 269086
rect 115764 269046 115916 269052
rect 115972 268921 116014 269124
rect 116164 269086 116316 269092
rect 116164 269052 116176 269086
rect 116304 269052 116316 269086
rect 116164 269046 116316 269052
rect 116372 268921 116414 269124
rect 116564 269086 116716 269092
rect 116564 269052 116576 269086
rect 116704 269052 116716 269086
rect 116564 269046 116716 269052
rect 116772 268921 116814 269124
rect 116964 269086 117116 269092
rect 116964 269052 116976 269086
rect 117104 269052 117116 269086
rect 116964 269046 117116 269052
rect 117172 268921 117214 269124
rect 117364 269086 117516 269092
rect 117364 269052 117376 269086
rect 117504 269052 117516 269086
rect 117364 269046 117516 269052
rect 117572 268921 117614 269124
rect 117764 269086 117916 269092
rect 117764 269052 117776 269086
rect 117904 269052 117916 269086
rect 117764 269046 117916 269052
rect 117972 268921 118014 269124
rect 118164 269086 118316 269092
rect 118164 269052 118176 269086
rect 118304 269052 118316 269086
rect 118164 269046 118316 269052
rect 118372 268921 118414 269124
rect 118564 269086 118716 269092
rect 118564 269052 118576 269086
rect 118704 269052 118716 269086
rect 118564 269046 118716 269052
rect 118772 268921 118814 269124
rect 120433 269130 120825 269136
rect 120433 269096 120445 269130
rect 120813 269096 120825 269130
rect 120433 269090 120825 269096
rect 121133 269130 121525 269136
rect 121133 269096 121145 269130
rect 121513 269096 121525 269130
rect 121133 269090 121525 269096
rect 112772 268888 118814 268921
rect 121991 268966 122023 269490
rect 122129 269374 122521 269380
rect 122129 269340 122141 269374
rect 122509 269340 122521 269374
rect 122129 269334 122521 269340
rect 122829 269374 123221 269380
rect 122829 269340 122841 269374
rect 123209 269340 123221 269374
rect 122829 269334 123221 269340
rect 122073 269281 122119 269293
rect 122073 269205 122079 269281
rect 122113 269205 122119 269281
rect 122073 269193 122119 269205
rect 122531 269281 122577 269293
rect 122531 269205 122537 269281
rect 122571 269205 122577 269281
rect 122531 269193 122577 269205
rect 122773 269281 122819 269293
rect 122773 269205 122779 269281
rect 122813 269205 122819 269281
rect 122773 269193 122819 269205
rect 123231 269281 123277 269293
rect 123231 269205 123237 269281
rect 123271 269205 123277 269281
rect 123231 269193 123277 269205
rect 122129 269146 122521 269152
rect 122129 269112 122141 269146
rect 122509 269112 122521 269146
rect 122129 269106 122521 269112
rect 122829 269146 123221 269152
rect 122829 269112 122841 269146
rect 123209 269112 123221 269146
rect 122829 269106 123221 269112
rect 123360 268966 123413 269638
rect 124192 269620 124204 269654
rect 124680 269620 124692 269654
rect 124192 269614 124692 269620
rect 124114 269592 124160 269604
rect 124114 269424 124120 269592
rect 124154 269424 124160 269592
rect 124114 269412 124160 269424
rect 124724 269592 124770 269608
rect 124724 269424 124730 269592
rect 124764 269424 124770 269592
rect 124724 269412 124770 269424
rect 124192 269396 124692 269402
rect 124192 269362 124204 269396
rect 124680 269362 124692 269396
rect 124192 269356 124692 269362
rect 121991 268908 123413 268966
rect 121991 268901 123412 268908
rect 114230 268883 117626 268888
rect 114230 268747 114322 268883
rect 117498 268747 117626 268883
rect 114230 268711 117626 268747
rect 125452 268342 125790 275158
rect 128055 268342 128452 275158
rect 125452 268022 128452 268342
rect 104286 266561 111587 266766
rect 104286 265524 104479 266561
rect 111335 265524 111587 266561
rect 104286 265368 111587 265524
<< via1 >>
rect 106140 282423 113415 283673
rect 102248 280847 103117 281654
rect 107422 279512 107721 279599
rect 108732 279512 109031 279599
rect 107381 279108 107553 279238
rect 102261 275681 103092 276478
rect 107015 277449 107487 277751
rect 107782 276842 107861 277125
rect 107978 276009 108049 276127
rect 109692 278009 109731 278872
rect 109731 278009 109744 278872
rect 109452 276623 109533 277299
rect 109687 276855 109731 277718
rect 109731 276855 109739 277718
rect 109918 276166 110180 276348
rect 109262 275859 109636 275949
rect 108227 275576 108353 275727
rect 114885 280226 114948 280294
rect 115257 280226 115320 280294
rect 114868 279813 114965 279861
rect 114965 279813 114966 279861
rect 114868 279809 114966 279813
rect 115239 279813 115240 279861
rect 115240 279813 115337 279861
rect 115239 279809 115337 279813
rect 114885 278560 114948 278628
rect 115257 278560 115320 278628
rect 119341 278715 119757 281145
rect 124552 280559 124902 280796
rect 120501 279564 120737 279656
rect 114868 278147 114965 278195
rect 114965 278147 114966 278195
rect 114868 278143 114966 278147
rect 115239 278147 115240 278195
rect 115240 278147 115337 278195
rect 115239 278143 115337 278147
rect 114885 276894 114948 276962
rect 115257 276894 115320 276962
rect 114868 276481 114965 276529
rect 114965 276481 114966 276529
rect 114868 276477 114966 276481
rect 115239 276481 115240 276529
rect 115240 276481 115337 276529
rect 115239 276477 115337 276481
rect 121605 277484 121657 279396
rect 121849 279275 122191 279887
rect 120958 276809 121013 277091
rect 114885 275228 114948 275296
rect 115257 275228 115320 275296
rect 114868 274815 114965 274863
rect 114965 274815 114966 274863
rect 114868 274811 114966 274815
rect 115239 274815 115240 274863
rect 115240 274815 115337 274863
rect 115239 274811 115337 274815
rect 102621 273772 105204 274070
rect 114885 273562 114948 273630
rect 115257 273562 115320 273630
rect 121822 276007 121912 276227
rect 122391 274783 122556 275289
rect 121823 273605 121913 273825
rect 114868 273149 114965 273197
rect 114965 273149 114966 273197
rect 114868 273145 114966 273149
rect 115239 273149 115240 273197
rect 115240 273149 115337 273197
rect 115239 273145 115337 273149
rect 122640 273395 122717 273451
rect 123785 273395 123862 273451
rect 107275 271829 107377 271953
rect 108641 272021 108841 272083
rect 107049 271327 107101 271473
rect 108445 271327 108497 271473
rect 106965 271115 107021 271313
rect 107049 270957 107101 271103
rect 108445 270957 108497 271103
rect 120958 272718 121013 273000
rect 114825 271918 115017 272012
rect 115017 271918 115527 272012
rect 114825 271817 115527 271918
rect 112267 270446 113449 270671
rect 121605 270428 121657 272340
rect 123380 272040 123463 272200
rect 124666 272845 124931 273042
rect 123962 270785 124063 271033
rect 123377 269673 123460 269833
rect 125790 268342 128055 275158
rect 104479 265524 111335 266561
<< metal2 >>
rect 105796 283673 113672 283895
rect 105796 282423 106140 283673
rect 113415 282423 113672 283673
rect 105796 282251 113672 282423
rect 102098 281654 103259 281810
rect 102098 280847 102248 281654
rect 103117 280847 103259 281654
rect 119257 281148 119845 281225
rect 121769 281148 122109 281149
rect 119257 281145 122109 281148
rect 102098 280720 103259 280847
rect 114322 281007 115149 281071
rect 114322 279876 114413 281007
rect 114865 280294 114970 280311
rect 114865 280226 114885 280294
rect 114948 280226 114970 280294
rect 114865 280204 114970 280226
rect 115069 280265 115149 281007
rect 115235 280294 115340 280311
rect 115235 280265 115257 280294
rect 115069 280226 115257 280265
rect 115320 280226 115340 280294
rect 115069 280213 115340 280226
rect 115235 280204 115340 280213
rect 114322 279861 115030 279876
rect 114322 279805 114868 279861
rect 114971 279805 115030 279861
rect 114322 279791 115030 279805
rect 115175 279861 115900 279876
rect 115175 279805 115234 279861
rect 115337 279805 115900 279861
rect 115175 279791 115900 279805
rect 107341 279599 107796 279642
rect 107341 279512 107422 279599
rect 107721 279512 107796 279599
rect 107341 279471 107796 279512
rect 108650 279599 109105 279641
rect 108650 279512 108732 279599
rect 109031 279554 109105 279599
rect 109031 279512 109575 279554
rect 108650 279491 109575 279512
rect 108650 279471 109576 279491
rect 107341 279238 107584 279471
rect 108978 279470 109576 279471
rect 107341 279108 107381 279238
rect 107553 279108 107584 279238
rect 107341 279074 107584 279108
rect 109441 278052 109576 279470
rect 109659 278872 109771 278903
rect 109659 278052 109692 278872
rect 109441 278009 109692 278052
rect 109744 278009 109771 278872
rect 114865 278628 114970 278645
rect 109441 277973 109771 278009
rect 114303 278560 114885 278628
rect 114948 278560 114970 278628
rect 114303 278543 114970 278560
rect 106957 277751 107553 277799
rect 106957 277449 107015 277751
rect 107487 277449 107553 277751
rect 109441 277755 109709 277973
rect 109441 277718 109771 277755
rect 109441 277695 109687 277718
rect 106957 277403 107553 277449
rect 109276 277299 109568 277341
rect 109276 277293 109452 277299
rect 107754 277125 107889 277153
rect 107754 276842 107782 277125
rect 107861 276842 107889 277125
rect 107754 276808 107889 276842
rect 102098 276478 103259 276621
rect 102098 275681 102261 276478
rect 103092 275681 103259 276478
rect 107789 276165 107889 276808
rect 109276 276695 109326 277293
rect 109276 276633 109452 276695
rect 109413 276623 109452 276633
rect 109533 276623 109568 277299
rect 109659 276855 109687 277695
rect 109739 276855 109771 277718
rect 109659 276825 109771 276855
rect 109413 276577 109568 276623
rect 114303 276544 114407 278543
rect 114865 278538 114970 278543
rect 115235 278632 115340 278645
rect 115788 278632 115900 279791
rect 115235 278628 115900 278632
rect 119257 278715 119341 281145
rect 119757 280610 122109 281145
rect 119757 278715 119845 280610
rect 121747 280609 122109 280610
rect 121899 279937 122109 280609
rect 124495 280796 124958 280846
rect 124495 280559 124552 280796
rect 124902 280559 124958 280796
rect 124495 280498 124958 280559
rect 121797 279887 122235 279937
rect 120433 279656 120825 279712
rect 120433 279564 120501 279656
rect 120737 279654 120825 279656
rect 120737 279564 121677 279654
rect 120433 279559 121677 279564
rect 120433 279510 120825 279559
rect 119257 278631 119845 278715
rect 121587 279396 121677 279559
rect 115235 278560 115257 278628
rect 115320 278560 115900 278628
rect 115235 278547 115900 278560
rect 115235 278538 115340 278547
rect 114843 278195 115030 278210
rect 114843 278139 114868 278195
rect 114971 278139 115030 278195
rect 114843 278125 115030 278139
rect 115175 278195 115362 278210
rect 115175 278139 115234 278195
rect 115337 278139 115362 278195
rect 115175 278125 115362 278139
rect 121587 277484 121605 279396
rect 121657 277814 121677 279396
rect 121797 279275 121849 279887
rect 122191 279275 122235 279887
rect 121797 279225 122235 279275
rect 121657 277718 121972 277814
rect 121657 277717 122169 277718
rect 121657 277504 122191 277717
rect 121657 277484 121677 277504
rect 121908 277503 122191 277504
rect 120953 277091 121018 277099
rect 114865 276962 114970 276979
rect 114865 276894 114885 276962
rect 114948 276894 114970 276962
rect 114865 276872 114970 276894
rect 115235 276962 115340 276979
rect 115235 276894 115257 276962
rect 115320 276894 115340 276962
rect 115235 276872 115340 276894
rect 120953 276809 120958 277091
rect 121013 276809 121018 277091
rect 114303 276529 115030 276544
rect 114303 276473 114868 276529
rect 114971 276473 115030 276529
rect 114303 276460 115030 276473
rect 114324 276459 115030 276460
rect 115175 276529 115900 276544
rect 115175 276473 115234 276529
rect 115337 276473 115900 276529
rect 115175 276459 115900 276473
rect 109383 276347 109700 276394
rect 109383 276165 109440 276347
rect 107789 276150 109440 276165
rect 109646 276165 109700 276347
rect 109824 276348 110271 276420
rect 109824 276166 109918 276348
rect 110180 276166 110271 276348
rect 109824 276165 110271 276166
rect 109646 276150 110271 276165
rect 107789 276127 110271 276150
rect 107789 276091 107978 276127
rect 107947 276009 107978 276091
rect 108049 276093 110271 276127
rect 108049 276091 109879 276093
rect 108049 276009 108079 276091
rect 107947 275970 108079 276009
rect 108280 275968 109712 275969
rect 108216 275949 109712 275968
rect 108216 275859 109262 275949
rect 109636 275859 109712 275949
rect 108216 275837 109712 275859
rect 108216 275765 108359 275837
rect 109193 275836 109712 275837
rect 102098 275531 103259 275681
rect 108187 275727 108393 275765
rect 108187 275576 108227 275727
rect 108353 275576 108393 275727
rect 108187 275522 108393 275576
rect 114865 275296 114970 275313
rect 114303 275228 114885 275296
rect 114948 275228 114970 275296
rect 114303 275211 114970 275228
rect 102557 274070 105283 274145
rect 102557 273772 102621 274070
rect 105204 273772 105283 274070
rect 102557 273716 105283 273772
rect 114303 273212 114407 275211
rect 114865 275206 114970 275211
rect 115235 275304 115340 275313
rect 115788 275304 115900 276459
rect 115235 275296 115900 275304
rect 115235 275228 115257 275296
rect 115320 275228 115900 275296
rect 115235 275219 115900 275228
rect 115235 275206 115340 275219
rect 114843 274863 115030 274878
rect 114843 274807 114868 274863
rect 114971 274807 115030 274863
rect 114843 274793 115030 274807
rect 115175 274863 115362 274878
rect 115175 274807 115234 274863
rect 115337 274807 115362 274863
rect 115175 274793 115362 274807
rect 114865 273632 114970 273647
rect 115235 273632 115340 273647
rect 114865 273630 115340 273632
rect 114865 273562 114885 273630
rect 114948 273562 115257 273630
rect 115320 273562 115340 273630
rect 114865 273554 115340 273562
rect 114865 273540 114970 273554
rect 115235 273540 115340 273554
rect 115209 273212 115899 273221
rect 114303 273197 115030 273212
rect 114303 273141 114868 273197
rect 114971 273141 115030 273197
rect 114303 273128 115030 273141
rect 114324 273127 115030 273128
rect 115175 273197 115899 273212
rect 115175 273141 115234 273197
rect 115337 273141 115899 273197
rect 115175 273127 115899 273141
rect 115209 273107 115899 273127
rect 104687 272547 108128 272685
rect 115759 272659 115899 273107
rect 120953 273000 121018 276809
rect 120953 272718 120958 273000
rect 121013 272718 121018 273000
rect 120953 272710 121018 272718
rect 115433 272645 115899 272659
rect 115433 272602 115898 272645
rect 104687 272454 108129 272547
rect 102092 271607 103253 271773
rect 102092 270822 102255 271607
rect 103070 271447 103253 271607
rect 104687 271447 104918 272454
rect 107985 272277 108129 272454
rect 107249 272207 108611 272277
rect 107249 271971 107351 272207
rect 108553 272113 108611 272207
rect 108553 272083 108841 272113
rect 108553 272021 108641 272083
rect 115433 272048 115559 272602
rect 121587 272340 121677 277484
rect 121801 276227 121931 276287
rect 121801 276007 121822 276227
rect 121912 276145 121931 276227
rect 121912 276007 121932 276145
rect 121801 275945 121932 276007
rect 121802 273825 121932 275945
rect 121802 273605 121823 273825
rect 121913 273605 121932 273825
rect 121802 273253 121932 273605
rect 122077 273466 122191 277503
rect 122326 275319 122757 275386
rect 122326 274780 122383 275319
rect 122718 274780 122757 275319
rect 122326 274706 122757 274780
rect 122602 273466 122755 273468
rect 122077 273451 122755 273466
rect 122077 273395 122640 273451
rect 122717 273449 122755 273451
rect 123747 273451 123900 273468
rect 123747 273449 123785 273451
rect 122717 273402 123785 273449
rect 122717 273395 122755 273402
rect 122077 273390 122755 273395
rect 122602 273371 122755 273390
rect 123747 273395 123785 273402
rect 123862 273395 123900 273451
rect 123747 273371 123900 273395
rect 121802 273151 123740 273253
rect 108553 271995 108841 272021
rect 114761 272012 115601 272048
rect 107249 271953 107401 271971
rect 107249 271829 107275 271953
rect 107377 271829 107401 271953
rect 107249 271807 107401 271829
rect 114761 271817 114825 272012
rect 115527 271817 115601 272012
rect 114761 271763 115601 271817
rect 103070 271216 104918 271447
rect 106951 271473 107141 271485
rect 106951 271327 107049 271473
rect 107101 271327 107141 271473
rect 106951 271315 107141 271327
rect 108405 271473 108507 271485
rect 108405 271327 108445 271473
rect 108497 271327 108507 271473
rect 108405 271315 108507 271327
rect 106951 271313 107095 271315
rect 103070 270822 103253 271216
rect 106951 271115 106965 271313
rect 107021 271115 107095 271313
rect 108451 271115 108507 271315
rect 106951 271103 107141 271115
rect 106951 270957 107049 271103
rect 107101 270957 107141 271103
rect 106951 270945 107141 270957
rect 108405 271103 108507 271115
rect 108405 270957 108445 271103
rect 108497 270957 108507 271103
rect 108405 270945 108507 270957
rect 102092 270683 103253 270822
rect 112194 270671 113508 270715
rect 112194 270446 112267 270671
rect 113449 270446 113508 270671
rect 112194 270399 113508 270446
rect 121587 270428 121605 272340
rect 121657 270428 121677 272340
rect 123362 272200 123476 272233
rect 123362 272040 123380 272200
rect 123463 272040 123476 272200
rect 123362 272007 123476 272040
rect 112198 267513 112378 270399
rect 121587 270345 121677 270428
rect 123381 269864 123456 272007
rect 123629 271620 123739 273151
rect 124813 273071 124957 280498
rect 124634 273042 124957 273071
rect 124634 272845 124666 273042
rect 124931 272849 124957 273042
rect 125452 275158 128452 275523
rect 124931 272845 124956 272849
rect 124634 272811 124956 272845
rect 123629 271526 124017 271620
rect 123629 271524 123739 271526
rect 123940 271093 124017 271526
rect 123931 271033 124081 271093
rect 123931 270785 123962 271033
rect 124063 270785 124081 271033
rect 123931 270717 124081 270785
rect 123360 269833 123474 269864
rect 123360 269673 123377 269833
rect 123460 269673 123474 269833
rect 123360 269638 123474 269673
rect 125452 268342 125790 275158
rect 128055 268342 128452 275158
rect 125452 268022 128452 268342
rect 112198 267463 116858 267513
rect 112198 267361 112243 267463
rect 116805 267361 116858 267463
rect 112198 267333 116858 267361
rect 104286 266561 111587 266766
rect 104286 265524 104479 266561
rect 111335 265524 111587 266561
rect 104286 265368 111587 265524
<< via2 >>
rect 106140 282423 113415 283673
rect 102248 280847 103117 281654
rect 114885 280226 114948 280294
rect 115257 280226 115320 280294
rect 114868 279809 114966 279861
rect 114966 279809 114971 279861
rect 114868 279805 114971 279809
rect 115234 279809 115239 279861
rect 115239 279809 115337 279861
rect 115234 279805 115337 279809
rect 114885 278560 114948 278628
rect 107015 277449 107487 277751
rect 102261 275681 103092 276478
rect 109326 276695 109452 277293
rect 109452 276695 109523 277293
rect 115257 278560 115320 278628
rect 114868 278143 114966 278195
rect 114966 278143 114971 278195
rect 114868 278139 114971 278143
rect 115234 278143 115239 278195
rect 115239 278143 115337 278195
rect 115234 278139 115337 278143
rect 114885 276894 114948 276962
rect 115257 276894 115320 276962
rect 114868 276477 114966 276529
rect 114966 276477 114971 276529
rect 114868 276473 114971 276477
rect 115234 276477 115239 276529
rect 115239 276477 115337 276529
rect 115234 276473 115337 276477
rect 109440 276150 109646 276347
rect 114885 275228 114948 275296
rect 102621 273772 105204 274070
rect 115257 275228 115320 275296
rect 114868 274811 114966 274863
rect 114966 274811 114971 274863
rect 114868 274807 114971 274811
rect 115234 274811 115239 274863
rect 115239 274811 115337 274863
rect 115234 274807 115337 274811
rect 114885 273562 114948 273630
rect 115257 273562 115320 273630
rect 114868 273145 114966 273197
rect 114966 273145 114971 273197
rect 114868 273141 114971 273145
rect 115234 273145 115239 273197
rect 115239 273145 115337 273197
rect 115234 273141 115337 273145
rect 102255 270822 103070 271607
rect 122383 275289 122718 275319
rect 122383 274783 122391 275289
rect 122391 274783 122556 275289
rect 122556 274783 122718 275289
rect 122383 274780 122718 274783
rect 125790 268342 128055 275158
rect 112243 267361 116805 267463
rect 104479 265524 111335 266561
<< metal3 >>
rect 572176 406600 582975 406686
rect 572176 406488 583606 406600
rect 572176 406300 582975 406488
rect 572176 374237 572562 406300
rect 154704 373851 572562 374237
rect 5373 337581 128286 337911
rect 344 337472 128286 337581
rect 5373 336821 128286 337472
rect 2990 294360 109888 295024
rect 342 294248 109888 294360
rect 2990 293144 109888 294248
rect 106790 283895 109888 293144
rect 105796 283673 113672 283895
rect 105796 282423 106140 283673
rect 113415 282423 113672 283673
rect 105796 282251 113672 282423
rect 127196 281912 128286 336821
rect 102098 281808 103259 281810
rect 6645 281654 103259 281808
rect 6645 280847 102248 281654
rect 103117 280847 103259 281654
rect 6645 280720 103259 280847
rect 127196 280822 128357 281912
rect 6645 280718 102170 280720
rect 6645 251338 7735 280718
rect 101936 280716 102170 280718
rect 114841 280294 114994 280329
rect 114303 280226 114885 280294
rect 114948 280226 114994 280294
rect 114303 280209 114994 280226
rect 106368 279497 109401 279505
rect 102586 279375 109401 279497
rect 102586 279266 106453 279375
rect 102586 279087 102817 279266
rect 107943 279238 109115 279266
rect 342 251226 7735 251338
rect 6645 251087 7735 251226
rect 31331 277997 103259 279087
rect 31331 124117 32421 277997
rect 106957 277751 107553 277799
rect 106957 277449 107015 277751
rect 107487 277449 107553 277751
rect 106957 277403 107553 277449
rect 102098 276620 103259 276621
rect 3945 123716 32421 124117
rect 326 123604 32421 123716
rect 3945 123027 32421 123604
rect 61553 276478 103259 276620
rect 61553 275681 102261 276478
rect 103092 275681 103259 276478
rect 107943 276214 107963 279238
rect 108027 276214 109115 279238
rect 109276 277341 109401 279375
rect 114303 278210 114407 280209
rect 114841 280178 114994 280209
rect 115211 280294 115364 280329
rect 115211 280226 115257 280294
rect 115320 280226 115364 280294
rect 115211 280178 115364 280226
rect 123842 279968 124731 280304
rect 127248 279968 127999 280822
rect 114843 279861 115030 279876
rect 114843 279805 114868 279861
rect 114971 279805 115030 279861
rect 114843 279791 115030 279805
rect 115175 279861 115362 279876
rect 115175 279805 115234 279861
rect 115337 279805 115362 279861
rect 115175 279791 115362 279805
rect 123842 279217 127999 279968
rect 123842 278876 124731 279217
rect 114841 278628 114994 278663
rect 114841 278560 114885 278628
rect 114948 278560 114994 278628
rect 114841 278512 114994 278560
rect 115211 278628 115364 278663
rect 115211 278560 115257 278628
rect 115320 278560 115364 278628
rect 115211 278512 115364 278560
rect 114303 278195 115030 278210
rect 114303 278139 114868 278195
rect 114971 278139 115030 278195
rect 114303 278126 115030 278139
rect 114324 278125 115030 278126
rect 115175 278195 115903 278210
rect 115175 278139 115234 278195
rect 115337 278139 115903 278195
rect 115175 278125 115903 278139
rect 109276 277293 109568 277341
rect 109276 276695 109326 277293
rect 109523 276695 109568 277293
rect 114841 276962 114994 276997
rect 109276 276633 109568 276695
rect 114303 276894 114885 276962
rect 114948 276894 114994 276962
rect 114303 276877 114994 276894
rect 107943 276186 109115 276214
rect 109383 276347 109700 276394
rect 109383 276150 109440 276347
rect 109646 276150 109700 276347
rect 109383 276091 109700 276150
rect 61553 275531 103259 275681
rect 61553 275530 102104 275531
rect 61553 80603 62643 275530
rect 114303 274878 114407 276877
rect 114841 276846 114994 276877
rect 115211 276972 115364 276997
rect 115791 276972 115903 278125
rect 124547 278165 124731 278876
rect 124547 277887 125086 278165
rect 115211 276962 115903 276972
rect 115211 276894 115257 276962
rect 115320 276894 115903 276962
rect 115211 276887 115903 276894
rect 115211 276846 115364 276887
rect 114843 276529 115030 276544
rect 114843 276473 114868 276529
rect 114971 276473 115030 276529
rect 114843 276459 115030 276473
rect 115175 276529 115362 276544
rect 115175 276473 115234 276529
rect 115337 276473 115362 276529
rect 115175 276459 115362 276473
rect 122326 275377 122757 275386
rect 124892 275377 125086 277887
rect 114841 275296 114994 275331
rect 114841 275228 114885 275296
rect 114948 275228 114994 275296
rect 114841 275180 114994 275228
rect 115211 275296 115364 275331
rect 115211 275228 115257 275296
rect 115320 275228 115364 275296
rect 115211 275180 115364 275228
rect 122326 275319 125086 275377
rect 114303 274863 115030 274878
rect 114303 274807 114868 274863
rect 114971 274807 115030 274863
rect 114303 274794 115030 274807
rect 114324 274793 115030 274794
rect 115175 274877 115362 274878
rect 115175 274863 115902 274877
rect 115175 274807 115234 274863
rect 115337 274807 115902 274863
rect 115175 274793 115902 274807
rect 115214 274792 115902 274793
rect 1853 80494 62643 80603
rect 342 80382 62643 80494
rect 1853 79513 62643 80382
rect 74033 274145 102558 274146
rect 74033 274070 105283 274145
rect 74033 273772 102621 274070
rect 105204 273772 105283 274070
rect 74033 273716 105283 273772
rect 1115 37272 4017 37406
rect 342 37245 4017 37272
rect 74033 37245 74463 273716
rect 114841 273630 114994 273665
rect 114841 273562 114885 273630
rect 114948 273562 114994 273630
rect 114841 273514 114994 273562
rect 115211 273635 115364 273665
rect 115790 273635 115902 274792
rect 122326 274780 122383 275319
rect 122718 275090 125086 275319
rect 125452 275158 128452 275523
rect 122718 274780 122757 275090
rect 122326 274706 122757 274780
rect 115211 273630 115902 273635
rect 115211 273562 115257 273630
rect 115320 273562 115902 273630
rect 115211 273550 115902 273562
rect 115211 273514 115364 273550
rect 114843 273197 115030 273212
rect 114843 273141 114868 273197
rect 114971 273141 115030 273197
rect 114843 273127 115030 273141
rect 115175 273197 115362 273212
rect 115175 273141 115234 273197
rect 115337 273141 115362 273197
rect 115175 273127 115362 273141
rect 342 37160 74463 37245
rect 1115 36815 74463 37160
rect 87083 271607 103253 271773
rect 87083 270822 102255 271607
rect 103070 270822 103253 271607
rect 87083 270683 103253 270822
rect 1115 36682 4017 36815
rect 87083 16181 88173 270683
rect 125452 268342 125790 275158
rect 128055 274476 128452 275158
rect 134328 274476 139500 350418
rect 128055 269304 139500 274476
rect 128055 268342 128452 269304
rect 125452 268022 128452 268342
rect 112198 267463 116858 267513
rect 112198 267361 112243 267463
rect 116805 267361 116858 267463
rect 112198 267333 116858 267361
rect 104286 266561 111587 266766
rect 104286 265524 104479 266561
rect 111335 265524 111587 266561
rect 104286 265368 111587 265524
rect 106618 236639 109716 265368
rect 115987 257334 116373 267333
rect 154704 257334 155090 373851
rect 115987 256948 155090 257334
rect 162337 364696 578379 366371
rect 162337 364584 581142 364696
rect 162337 363273 578379 364584
rect 162337 236639 165435 363273
rect 581030 360178 581142 364584
rect 581030 360066 583606 360178
rect 106618 233541 165435 236639
rect 1455 15850 88173 16181
rect 342 15738 88173 15850
rect 1455 15091 88173 15738
<< via3 >>
rect 107015 277449 107487 277751
rect 107963 276214 108027 279238
rect 109440 276150 109646 276347
<< mimcap >>
rect 108275 279186 109075 279226
rect 108275 276266 108315 279186
rect 109035 276266 109075 279186
rect 108275 276226 109075 276266
<< mimcapcontact >>
rect 108315 276266 109035 279186
<< metal4 >>
rect 107947 279238 108043 279254
rect 106957 277751 107553 277799
rect 106957 277449 107015 277751
rect 107487 277737 107553 277751
rect 107947 277737 107963 279238
rect 107487 277477 107963 277737
rect 107487 277449 107553 277477
rect 106957 277403 107553 277449
rect 107947 276214 107963 277477
rect 108027 276214 108043 279238
rect 108314 279186 109036 279187
rect 108314 276266 108315 279186
rect 109035 276394 109036 279186
rect 109035 276347 109700 276394
rect 109035 276266 109440 276347
rect 108314 276265 109440 276266
rect 107947 276198 108043 276214
rect 109383 276150 109440 276265
rect 109646 276150 109700 276347
rect 109383 276091 109700 276150
<< labels >>
flabel metal3 10028 336906 11894 337768 0 FreeSans 8000 0 0 0 gpio_noesd[11]
port 0 nsew
flabel metal3 9412 293530 11278 294392 0 FreeSans 8000 0 0 0 gpio_noesd[12]
port 1 nsew
flabel metal3 6760 251254 7466 251912 0 FreeSans 8000 0 0 0 gpio_noesd[13]
port 2 nsew
flabel metal3 7748 123292 8454 123950 0 FreeSans 8000 0 0 0 gpio_noesd[14]
port 3 nsew
flabel metal3 7280 79630 7986 80288 0 FreeSans 8000 0 0 0 gpio_noesd[15]
port 4 nsew
flabel metal3 6896 36870 8062 37110 0 FreeSans 8000 0 0 0 gpio_noesd[16]
port 5 nsew
flabel metal3 6686 15490 7852 15730 0 FreeSans 8000 0 0 0 gpio_noesd[17]
port 6 nsew
flabel metal3 573308 364318 574122 364838 0 FreeSans 8000 0 0 0 gpio_noesd[2]
port 7 nsew
flabel metal3 575802 406322 576204 406584 0 FreeSans 8000 0 0 0 gpio_noesd[3]
port 8 nsew
flabel metal3 135612 346104 138678 348766 0 FreeSans 12800 0 0 0 vssa1
port 9 nsew
flabel metal2 112229 267697 112349 267811 0 FreeSans 3200 90 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_out
flabel metal1 111201 267695 111321 267809 0 FreeSans 3200 90 0 0 pmu_circuits_top_level_0/pmu_circuits_0.dd_02
flabel metal2 106605 272511 106725 272625 0 FreeSans 3200 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.vref
flabel metal1 106117 277553 106237 277667 0 FreeSans 3200 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_out
flabel metal1 105863 278241 105937 278329 0 FreeSans 3200 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_vs
flabel metal3 105859 279345 105933 279433 0 FreeSans 3200 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_vb
flabel metal1 105821 281133 105895 281221 0 FreeSans 3200 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_iref
flabel metal1 106163 282527 106237 282615 0 FreeSans 3200 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.dd_01
flabel locali 125137 281485 125329 281667 0 FreeSans 3200 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ss
flabel metal3 125259 279535 125451 279717 0 FreeSans 3200 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref
flabel metal2 108523 272221 108591 272269 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.vref01_0.VREF
flabel metal1 108587 270871 108655 270919 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.vref01_0.DD
flabel locali 106809 271879 106877 271927 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.vref01_0.SS
flabel locali 118007 272352 118355 272604 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.SS
flabel metal1 113347 272304 113553 272494 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.DD
flabel space 112715 270440 112921 270630 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.OUT
flabel metal1 112489 270487 112617 270591 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.ring_100mV_buffer_0.OUT
flabel metal2 114788 271797 114916 271901 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.ring_100mV_buffer_0.IN
flabel viali 113883 271822 114011 271926 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.ring_100mV_buffer_0.DD
flabel locali 119001 272134 119129 272238 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.ring_100mV_buffer_0.SS
rlabel metal1 114297 279009 114372 279073 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_9.IN
rlabel locali 113345 277680 113420 277744 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_9.SS
rlabel locali 114959 277764 114997 277798 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_9.DD
rlabel metal1 112782 277799 112826 277838 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_9.OUT
rlabel metal1 115833 279009 115908 279073 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_8.IN
rlabel locali 116785 277680 116860 277744 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_8.SS
rlabel locali 115208 277764 115246 277798 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_8.DD
rlabel metal1 117379 277799 117423 277838 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_8.OUT
rlabel metal1 114297 277343 114372 277407 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_7.IN
rlabel locali 113345 276014 113420 276078 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_7.SS
rlabel locali 114959 276098 114997 276132 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_7.DD
rlabel metal1 112782 276133 112826 276172 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT
rlabel metal1 115833 277343 115908 277407 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN
rlabel locali 116785 276014 116860 276078 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_6.SS
rlabel locali 115208 276098 115246 276132 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_6.DD
rlabel metal1 117379 276133 117423 276172 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_6.OUT
rlabel metal1 114297 275677 114372 275741 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_5.IN
rlabel locali 113345 274348 113420 274412 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_5.SS
rlabel locali 114959 274432 114997 274466 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_5.DD
rlabel metal1 112782 274467 112826 274506 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT
rlabel metal1 115833 275677 115908 275741 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN
rlabel locali 116785 274348 116860 274412 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_4.SS
rlabel locali 115208 274432 115246 274466 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_4.DD
rlabel metal1 117379 274467 117423 274506 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_4.OUT
rlabel metal1 115833 274011 115908 274075 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_3.IN
rlabel locali 116785 272682 116860 272746 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_3.SS
rlabel locali 115208 272766 115246 272800 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_3.DD
rlabel metal1 117379 272801 117423 272840 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT
rlabel metal1 114297 274011 114372 274075 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN
rlabel locali 113345 272682 113420 272746 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_2.SS
rlabel locali 114959 272766 114997 272800 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_2.DD
rlabel metal1 112782 272801 112826 272840 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT
rlabel metal1 115833 280675 115908 280739 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_1.IN
rlabel locali 116785 279346 116860 279410 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_1.SS
rlabel locali 115208 279430 115246 279464 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_1.DD
rlabel metal1 117379 279465 117423 279504 7 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT
rlabel metal1 114297 280675 114372 280739 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN
rlabel locali 113345 279346 113420 279410 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_0.SS
rlabel locali 114959 279430 114997 279464 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_0.DD
rlabel metal1 112782 279465 112826 279504 3 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT
flabel metal1 108183 280591 108259 280679 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_0.Iref
flabel locali 109921 279361 109997 279449 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_0.SS
flabel metal3 106173 279327 106347 279459 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_0.VB
flabel metal1 106071 278255 106121 278309 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_0.VS
flabel metal1 106327 277543 106527 277719 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_0.OUT
flabel metal1 106143 274775 106235 274891 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_0.DD
flabel metal2 120471 280709 120701 280913 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.DD
flabel metal3 124171 279421 124401 279625 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.IREF
flabel locali 123893 268977 124041 269141 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.SS
flabel locali 122378 278528 122456 278606 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_vref_0.DD
flabel locali 122060 276558 122134 276644 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_vref_0.SS
flabel metal1 124468 276546 124542 276632 0 FreeSans 1600 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_vref_0.VREF
rlabel metal2 121796 277545 121931 277755 1 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Ip2
rlabel metal1 121951 274874 122001 274947 1 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Iref
rlabel metal1 123719 270947 123769 271020 1 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Vg
rlabel metal2 123405 269727 123455 269800 1 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Ip1
rlabel locali 124373 269012 124499 269117 1 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.SS
rlabel locali 121944 279849 122032 279923 1 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.DD
rlabel metal1 124871 273456 124913 273514 3 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg
rlabel metal1 123437 273648 123479 273706 3 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1
rlabel metal1 123851 273648 123893 273706 3 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2
rlabel locali 124019 274734 124061 274792 3 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.SS
rlabel metal1 124223 274754 124265 274812 3 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT
<< end >>

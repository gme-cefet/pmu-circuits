magic
tech sky130A
magscale 1 2
timestamp 1698328593
<< error_s >>
rect 12527 -8940 12530 -8906
rect 12561 -8974 12564 -8872
<< nwell >>
rect 9004 -5155 12217 -3862
rect 11083 -8443 12754 -7099
<< psubdiff >>
rect 8663 -3804 8720 -3712
rect 12773 -3804 12913 -3712
rect 8663 -3854 8742 -3804
rect 12827 -3820 12913 -3804
rect 8663 -5733 8742 -5241
rect 8700 -8726 8834 -8355
rect 8574 -8810 8659 -8726
rect 12717 -8810 12827 -8726
rect 8574 -8883 8656 -8810
rect 8574 -10146 8656 -10047
rect 12680 -8901 12827 -8810
rect 12762 -10065 12827 -8901
rect 12680 -10146 12827 -10065
rect 8574 -10230 8659 -10146
rect 12717 -10226 12827 -10146
rect 12717 -10230 12913 -10226
rect 12740 -10250 12913 -10230
<< nsubdiff >>
rect 9040 -3932 9100 -3898
rect 12121 -3932 12181 -3898
rect 9040 -3958 9074 -3932
rect 9040 -5085 9074 -5059
rect 12147 -3958 12181 -3932
rect 12147 -5085 12181 -5059
rect 9040 -5119 9100 -5085
rect 12121 -5119 12181 -5085
rect 11119 -7169 11179 -7135
rect 12658 -7169 12718 -7135
rect 11119 -7195 11153 -7169
rect 11119 -8373 11153 -8347
rect 12684 -7195 12718 -7169
rect 12684 -8373 12718 -8347
rect 11119 -8407 11179 -8373
rect 12658 -8407 12718 -8373
<< psubdiffcont >>
rect 8720 -3804 12773 -3712
rect 8663 -5241 8742 -3854
rect 8659 -8810 12717 -8726
rect 8574 -10047 8656 -8883
rect 12680 -10065 12762 -8901
rect 8659 -10230 12717 -10146
rect 12827 -10226 12913 -3820
<< nsubdiffcont >>
rect 9100 -3932 12121 -3898
rect 9040 -5059 9074 -3958
rect 12147 -5059 12181 -3958
rect 9100 -5119 12121 -5085
rect 11179 -7169 12658 -7135
rect 11119 -8347 11153 -7195
rect 12684 -8347 12718 -7195
rect 11179 -8407 12658 -8373
<< locali >>
rect 8663 -3804 8720 -3712
rect 12773 -3804 12913 -3712
rect 8663 -3854 8742 -3804
rect 12827 -3820 12913 -3804
rect 9040 -3932 9100 -3898
rect 12121 -3916 12181 -3898
rect 12121 -3932 12593 -3916
rect 9040 -3958 12593 -3932
rect 9074 -4067 12147 -3958
rect 9074 -4251 9195 -4067
rect 9254 -4071 12147 -4067
rect 9254 -4074 11940 -4071
rect 9074 -4732 9191 -4251
rect 11996 -4264 12147 -4071
rect 12013 -4726 12147 -4264
rect 9074 -5059 9194 -4732
rect 9040 -5085 9194 -5059
rect 9309 -5085 9389 -4927
rect 11812 -5085 11892 -4924
rect 12000 -5059 12147 -4726
rect 12181 -4038 12593 -3958
rect 12181 -5059 12338 -4038
rect 12000 -5085 12338 -5059
rect 9040 -5119 9100 -5085
rect 12121 -5119 12338 -5085
rect 8663 -5738 8742 -5241
rect 8575 -5740 8742 -5738
rect 11902 -5475 12338 -5119
rect 12512 -5475 12593 -4038
rect 11902 -5588 12593 -5475
rect 8575 -8356 8683 -5740
rect 11902 -6124 12168 -5588
rect 11902 -6131 12130 -6124
rect 11754 -6246 12038 -6140
rect 11757 -6974 11985 -6909
rect 11757 -7135 11789 -6974
rect 11946 -7135 11985 -6974
rect 11119 -7169 11179 -7135
rect 12658 -7169 12718 -7135
rect 11119 -7195 11153 -7169
rect 11650 -7253 11789 -7169
rect 11946 -7253 12125 -7169
rect 11650 -7311 12125 -7253
rect 12684 -7195 12718 -7169
rect 11212 -8196 11258 -7342
rect 12566 -8196 12612 -7342
rect 8575 -8726 9251 -8356
rect 11119 -8373 11153 -8347
rect 12684 -8373 12718 -8347
rect 11119 -8407 11179 -8373
rect 12658 -8407 12718 -8373
rect 8574 -8810 8659 -8726
rect 12717 -8734 12762 -8726
rect 12717 -8810 12827 -8734
rect 8574 -8883 8905 -8810
rect 8656 -8923 8905 -8883
rect 9198 -8906 12130 -8872
rect 8656 -8932 8880 -8923
rect 8656 -9319 8758 -8932
rect 8930 -8974 8976 -8906
rect 12352 -8974 12398 -8906
rect 12424 -8923 12506 -8810
rect 12561 -8901 12827 -8810
rect 8656 -9713 8777 -9319
rect 8656 -10036 8758 -9713
rect 8656 -10047 8799 -10036
rect 8574 -10061 8799 -10047
rect 8825 -10061 8907 -10050
rect 8574 -10146 8907 -10061
rect 9107 -10146 9152 -8974
rect 9507 -10146 9552 -8974
rect 9907 -10146 9952 -8974
rect 10307 -10146 10352 -8974
rect 10976 -10146 11021 -8974
rect 11376 -10146 11421 -8974
rect 11776 -10146 11821 -8974
rect 12176 -10146 12221 -8974
rect 12561 -9934 12680 -8901
rect 12542 -10036 12680 -9934
rect 12473 -10046 12680 -10036
rect 12422 -10065 12680 -10046
rect 12762 -10065 12827 -8901
rect 12422 -10146 12827 -10065
rect 8574 -10230 8659 -10146
rect 12717 -10226 12827 -10146
rect 12717 -10230 12913 -10226
rect 12666 -10249 12913 -10230
<< viali >>
rect 12338 -5475 12512 -4038
rect 11789 -7135 11946 -6974
rect 11789 -7169 11946 -7135
rect 11789 -7253 11946 -7169
<< metal1 >>
rect 12265 -3916 12787 -3841
rect 12264 -4038 12787 -3916
rect 10005 -4578 10193 -4444
rect 10505 -4578 10693 -4444
rect 11005 -4578 11193 -4444
rect 10506 -4761 10686 -4707
rect 10506 -4894 10534 -4761
rect 10436 -4912 10534 -4894
rect 10660 -4894 10686 -4761
rect 10660 -4912 10758 -4894
rect 9820 -5017 9880 -4916
rect 10436 -4950 10758 -4912
rect 11320 -5017 11380 -4916
rect 9175 -5044 9694 -5021
rect 9175 -5134 9251 -5044
rect 9625 -5134 9694 -5044
rect 9820 -5067 11380 -5017
rect 9175 -5154 9694 -5134
rect 8616 -5351 9063 -5278
rect 8616 -5533 8707 -5351
rect 8969 -5533 9063 -5351
rect 8616 -5605 9063 -5533
rect 8631 -5902 8738 -5605
rect 8828 -5808 9474 -5762
rect 8828 -5824 9354 -5808
rect 8631 -7245 8772 -5902
rect 9116 -6040 9228 -6010
rect 9116 -6903 9148 -6040
rect 9200 -6903 9228 -6040
rect 9116 -6940 9228 -6903
rect 9318 -6484 9354 -5824
rect 9435 -6484 9474 -5808
rect 9318 -6526 9474 -6484
rect 9318 -7018 9370 -6526
rect 8828 -7080 9370 -7018
rect 8722 -8196 8772 -7245
rect 9116 -7194 9228 -7158
rect 9116 -8057 9143 -7194
rect 9195 -8057 9228 -7194
rect 9116 -8088 9228 -8057
rect 9318 -8274 9370 -7080
rect 8828 -8336 9370 -8274
rect 9596 -8533 9691 -5154
rect 10808 -5194 10940 -5067
rect 10808 -5312 10838 -5194
rect 10909 -5312 10940 -5194
rect 10808 -5350 10940 -5312
rect 12264 -5475 12338 -4038
rect 12512 -4522 12787 -4038
rect 12512 -5475 12593 -4522
rect 12264 -5588 12593 -5475
rect 10998 -6027 12483 -5993
rect 10998 -6310 11026 -6027
rect 11105 -6040 12483 -6027
rect 11105 -6287 11133 -6040
rect 11105 -6310 11292 -6287
rect 10998 -6343 11292 -6310
rect 12437 -6345 12483 -6040
rect 11806 -6588 11928 -6374
rect 11334 -6592 11930 -6588
rect 12127 -6592 12718 -6582
rect 11334 -6634 12718 -6592
rect 11334 -6936 11400 -6634
rect 11872 -6812 12718 -6634
rect 11872 -6909 11930 -6812
rect 11872 -6936 11985 -6909
rect 11334 -6974 11985 -6936
rect 11334 -6984 11789 -6974
rect 11757 -7223 11789 -6984
rect 11091 -7253 11789 -7223
rect 11946 -7223 11985 -6974
rect 12127 -7010 12718 -6812
rect 11946 -7253 12519 -7223
rect 11091 -7290 12519 -7253
rect 11091 -7823 11178 -7290
rect 12590 -7564 12821 -7364
rect 11305 -7715 12739 -7648
rect 11091 -7890 12519 -7823
rect 12652 -8248 12739 -7715
rect 11305 -8250 12739 -8248
rect 11303 -8293 12739 -8250
rect 11303 -8423 11334 -8293
rect 11506 -8315 12739 -8293
rect 11506 -8423 11547 -8315
rect 11303 -8443 11547 -8423
rect 9382 -8586 11946 -8533
rect 9382 -9998 9437 -8586
rect 9782 -8697 11546 -8656
rect 9782 -8784 9856 -8697
rect 10155 -8704 11166 -8697
rect 10155 -8784 10237 -8704
rect 9782 -8826 10237 -8784
rect 9782 -9998 9837 -8826
rect 10182 -9998 10237 -8826
rect 11091 -8784 11166 -8704
rect 11465 -8784 11546 -8697
rect 11091 -8827 11546 -8784
rect 10582 -9998 10746 -8978
rect 11091 -9998 11146 -8827
rect 11491 -9998 11546 -8827
rect 11891 -9998 11946 -8586
rect 10632 -10064 10691 -9998
rect 9202 -10134 12126 -10064
rect 10592 -10258 10741 -10134
<< via1 >>
rect 10534 -4912 10660 -4761
rect 9251 -5134 9625 -5044
rect 8707 -5533 8969 -5351
rect 9148 -6903 9200 -6040
rect 9354 -6484 9435 -5808
rect 9143 -8057 9195 -7194
rect 10838 -5312 10909 -5194
rect 11026 -6310 11105 -6027
rect 11400 -6936 11872 -6634
rect 11334 -8423 11506 -8293
rect 9856 -8784 10155 -8697
rect 11166 -8784 11465 -8697
<< metal2 >>
rect 10494 -4761 10700 -4707
rect 10494 -4912 10534 -4761
rect 10660 -4912 10700 -4761
rect 10494 -4950 10700 -4912
rect 9175 -5022 9694 -5021
rect 10528 -5022 10671 -4950
rect 9175 -5044 10671 -5022
rect 9175 -5134 9251 -5044
rect 9625 -5134 10671 -5044
rect 9175 -5153 10671 -5134
rect 9175 -5154 10607 -5153
rect 10808 -5194 10940 -5155
rect 10808 -5276 10838 -5194
rect 9008 -5278 10838 -5276
rect 8616 -5312 10838 -5278
rect 10909 -5276 10940 -5194
rect 10909 -5312 11098 -5276
rect 8616 -5335 11098 -5312
rect 8616 -5350 9241 -5335
rect 8616 -5351 9063 -5350
rect 8616 -5533 8707 -5351
rect 8969 -5533 9063 -5351
rect 8616 -5605 9063 -5533
rect 9187 -5532 9241 -5350
rect 9447 -5350 11098 -5335
rect 9447 -5532 9504 -5350
rect 9187 -5579 9504 -5532
rect 9319 -5808 9474 -5762
rect 9116 -6040 9228 -6010
rect 9116 -6903 9148 -6040
rect 9200 -6880 9228 -6040
rect 9319 -6484 9354 -5808
rect 9435 -5818 9474 -5808
rect 9435 -5880 9611 -5818
rect 9561 -6478 9611 -5880
rect 10998 -5993 11098 -5350
rect 10998 -6027 11133 -5993
rect 10998 -6310 11026 -6027
rect 11105 -6310 11133 -6027
rect 10998 -6338 11133 -6310
rect 9435 -6484 9611 -6478
rect 9319 -6526 9611 -6484
rect 11334 -6634 11930 -6588
rect 9200 -6903 9446 -6880
rect 9116 -6940 9446 -6903
rect 9178 -7158 9446 -6940
rect 11334 -6936 11400 -6634
rect 11872 -6936 11930 -6634
rect 11334 -6984 11930 -6936
rect 9116 -7194 9446 -7158
rect 9116 -8057 9143 -7194
rect 9195 -7237 9446 -7194
rect 9195 -8057 9228 -7237
rect 9116 -8088 9228 -8057
rect 9311 -8655 9446 -7237
rect 11303 -8293 11546 -8259
rect 11303 -8423 11334 -8293
rect 11506 -8423 11546 -8293
rect 9311 -8656 9909 -8655
rect 11303 -8656 11546 -8423
rect 9311 -8676 10237 -8656
rect 9312 -8697 10237 -8676
rect 9312 -8739 9856 -8697
rect 9782 -8784 9856 -8739
rect 10155 -8784 10237 -8697
rect 9782 -8826 10237 -8784
rect 11091 -8697 11546 -8656
rect 11091 -8784 11166 -8697
rect 11465 -8784 11546 -8697
rect 11091 -8827 11546 -8784
<< via2 >>
rect 9241 -5532 9447 -5335
rect 9364 -6478 9435 -5880
rect 9435 -6478 9561 -5880
rect 11400 -6936 11872 -6634
<< metal3 >>
rect 9187 -5335 9504 -5276
rect 9187 -5532 9241 -5335
rect 9447 -5532 9504 -5335
rect 9187 -5579 9504 -5532
rect 9319 -5880 9611 -5818
rect 9319 -6478 9364 -5880
rect 9561 -6478 9611 -5880
rect 9319 -6526 9611 -6478
rect 9486 -8560 9611 -6526
rect 11334 -6634 11930 -6588
rect 11334 -6936 11400 -6634
rect 11872 -6936 11930 -6634
rect 11334 -6984 11930 -6936
rect 12434 -8560 12913 -8451
rect 9486 -8682 12913 -8560
rect 9486 -8690 12519 -8682
<< via3 >>
rect 9241 -5532 9447 -5335
rect 11400 -6936 11872 -6634
<< metal4 >>
rect 9187 -5335 9504 -5276
rect 9187 -5532 9241 -5335
rect 9447 -5450 9504 -5335
rect 9447 -5532 10120 -5450
rect 9187 -5579 10120 -5532
rect 11334 -6634 11930 -6588
rect 11334 -6662 11400 -6634
rect 10882 -6922 11400 -6662
rect 11334 -6936 11400 -6922
rect 11872 -6936 11930 -6634
rect 11334 -6984 11930 -6936
use sky130_fd_pr__cap_mim_m3_1_4FSB7X  sky130_fd_pr__cap_mim_m3_1_4FSB7X_0
timestamp 1696350080
transform 1 0 10358 0 1 -6911
box -586 -1540 586 1540
use sky130_fd_pr__nfet_01v8_lvt_5VYM7K  sky130_fd_pr__nfet_01v8_lvt_5VYM7K_0
timestamp 1696344833
transform 1 0 10864 0 1 -9488
box -124 -598 124 598
use sky130_fd_pr__nfet_01v8_lvt_5VYM7K  sky130_fd_pr__nfet_01v8_lvt_5VYM7K_1
timestamp 1696344833
transform 1 0 8864 0 1 -9488
box -124 -598 124 598
use sky130_fd_pr__nfet_01v8_lvt_5VYM7K  sky130_fd_pr__nfet_01v8_lvt_5VYM7K_2
timestamp 1696344833
transform 1 0 9264 0 1 -9488
box -124 -598 124 598
use sky130_fd_pr__nfet_01v8_lvt_5VYM7K  sky130_fd_pr__nfet_01v8_lvt_5VYM7K_3
timestamp 1696344833
transform 1 0 9664 0 1 -9488
box -124 -598 124 598
use sky130_fd_pr__nfet_01v8_lvt_5VYM7K  sky130_fd_pr__nfet_01v8_lvt_5VYM7K_4
timestamp 1696344833
transform 1 0 10064 0 1 -9488
box -124 -598 124 598
use sky130_fd_pr__nfet_01v8_lvt_5VYM7K  sky130_fd_pr__nfet_01v8_lvt_5VYM7K_5
timestamp 1696344833
transform 1 0 10464 0 1 -9488
box -124 -598 124 598
use sky130_fd_pr__nfet_01v8_lvt_5VYM7K  sky130_fd_pr__nfet_01v8_lvt_5VYM7K_6
timestamp 1696344833
transform 1 0 11664 0 1 -9488
box -124 -598 124 598
use sky130_fd_pr__nfet_01v8_lvt_5VYM7K  sky130_fd_pr__nfet_01v8_lvt_5VYM7K_7
timestamp 1696344833
transform 1 0 11264 0 1 -9488
box -124 -598 124 598
use sky130_fd_pr__nfet_01v8_lvt_5VYM7K  sky130_fd_pr__nfet_01v8_lvt_5VYM7K_8
timestamp 1696344833
transform 1 0 12464 0 1 -9488
box -124 -598 124 598
use sky130_fd_pr__nfet_01v8_lvt_5VYM7K  sky130_fd_pr__nfet_01v8_lvt_5VYM7K_9
timestamp 1696344833
transform 1 0 12064 0 1 -9488
box -124 -598 124 598
use sky130_fd_pr__nfet_01v8_lvt_W6ELF5  sky130_fd_pr__nfet_01v8_lvt_W6ELF5_0
timestamp 1696345916
transform 1 0 8967 0 1 -7049
box -339 -1357 339 1357
use sky130_fd_pr__pfet_01v8_lvt_8D4JM4  sky130_fd_pr__pfet_01v8_lvt_8D4JM4_0
timestamp 1696346853
transform 0 1 11912 -1 0 -7469
box -221 -707 221 707
use sky130_fd_pr__pfet_01v8_lvt_8D4JM4  sky130_fd_pr__pfet_01v8_lvt_8D4JM4_1
timestamp 1696346853
transform 0 1 11912 -1 0 -8069
box -221 -707 221 707
use sky130_fd_pr__pfet_01v8_lvt_EFQJD4  sky130_fd_pr__pfet_01v8_lvt_EFQJD4_0
timestamp 1696346853
transform 0 1 11879 -1 0 -6312
box -233 -736 233 736
use sky130_fd_pr__pfet_01v8_TRB9BZ  sky130_fd_pr__pfet_01v8_TRB9BZ_0
timestamp 1696340207
transform 0 1 11847 -1 0 -4509
box -483 -189 483 189
use sky130_fd_pr__pfet_01v8_TRB9BZ  sky130_fd_pr__pfet_01v8_TRB9BZ_1
timestamp 1696340207
transform 0 1 9347 -1 0 -4509
box -483 -189 483 189
use sky130_fd_pr__pfet_01v8_TRB9BZ  sky130_fd_pr__pfet_01v8_TRB9BZ_2
timestamp 1696340207
transform 0 1 9847 -1 0 -4509
box -483 -189 483 189
use sky130_fd_pr__pfet_01v8_TRB9BZ  sky130_fd_pr__pfet_01v8_TRB9BZ_3
timestamp 1696340207
transform 0 1 10347 -1 0 -4509
box -483 -189 483 189
use sky130_fd_pr__pfet_01v8_TRB9BZ  sky130_fd_pr__pfet_01v8_TRB9BZ_4
timestamp 1696340207
transform 0 1 10847 -1 0 -4509
box -483 -189 483 189
use sky130_fd_pr__pfet_01v8_TRB9BZ  sky130_fd_pr__pfet_01v8_TRB9BZ_5
timestamp 1696340207
transform 0 1 11347 -1 0 -4509
box -483 -189 483 189
<< labels >>
flabel metal1 10628 -9864 10704 -9776 0 FreeSans 1600 0 0 0 Iref
port 0 nsew
flabel locali 8890 -8634 8966 -8546 0 FreeSans 1600 0 0 0 SS
port 1 nsew
flabel metal3 12540 -8644 12714 -8512 0 FreeSans 1600 0 0 0 VB
port 2 nsew
flabel metal1 12766 -7494 12816 -7440 0 FreeSans 1600 0 0 0 VS
port 3 nsew
flabel metal1 12360 -6904 12560 -6728 0 FreeSans 1600 0 0 0 OUT
port 4 nsew
flabel metal1 12652 -4076 12744 -3960 0 FreeSans 1600 0 0 0 DD
port 5 nsew
<< end >>
